VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1429.100 2924.800 1430.300 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.650 3517.600 2229.210 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.810 3517.600 1905.370 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 3517.600 1581.530 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.290 3517.600 933.850 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.450 3517.600 610.010 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 3517.600 286.170 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3471.140 2.400 3472.340 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3212.740 2.400 3213.940 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2954.340 2.400 2955.540 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.940 2924.800 1694.140 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2695.940 2.400 2697.140 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2437.540 2.400 2438.740 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2179.140 2.400 2180.340 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1920.740 2.400 1921.940 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1662.340 2.400 1663.540 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1403.940 2.400 1405.140 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1145.540 2.400 1146.740 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 887.140 2.400 888.340 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 628.740 2.400 629.940 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1956.780 2924.800 1957.980 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2220.620 2924.800 2221.820 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2484.460 2924.800 2485.660 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2748.300 2924.800 2749.500 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3012.140 2924.800 3013.340 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3275.980 2924.800 3277.180 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.330 3517.600 2876.890 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2552.490 3517.600 2553.050 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 43.940 2924.800 45.140 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2286.580 2924.800 2287.780 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2550.420 2924.800 2551.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2814.260 2924.800 2815.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.100 2924.800 3079.300 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3341.940 2924.800 3343.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2795.370 3517.600 2795.930 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.530 3517.600 2472.090 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.690 3517.600 2148.250 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.850 3517.600 1824.410 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.010 3517.600 1500.570 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 241.820 2924.800 243.020 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.170 3517.600 1176.730 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.330 3517.600 852.890 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 3517.600 529.050 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 3517.600 205.210 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3148.140 2.400 3149.340 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2889.740 2.400 2890.940 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2631.340 2.400 2632.540 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2372.940 2.400 2374.140 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2114.540 2.400 2115.740 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.700 2924.800 440.900 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1597.740 2.400 1598.940 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1339.340 2.400 1340.540 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1080.940 2.400 1082.140 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 822.540 2.400 823.740 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 564.140 2.400 565.340 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 370.340 2.400 371.540 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 176.540 2.400 177.740 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 637.580 2924.800 638.780 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 835.460 2924.800 836.660 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1033.340 2924.800 1034.540 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1231.220 2924.800 1232.420 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2022.740 2924.800 2023.940 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 175.860 2924.800 177.060 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2418.500 2924.800 2419.700 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2682.340 2924.800 2683.540 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2946.180 2924.800 2947.380 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3210.020 2924.800 3211.220 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3473.860 2924.800 3475.060 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2633.450 3517.600 2634.010 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.610 3517.600 2310.170 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.770 3517.600 1986.330 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 3517.600 1662.490 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 373.740 2924.800 374.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.250 3517.600 1014.810 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.410 3517.600 690.970 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.570 3517.600 367.130 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.730 3517.600 43.290 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3277.340 2.400 3278.540 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3018.940 2.400 3020.140 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2760.540 2.400 2761.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2502.140 2.400 2503.340 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2243.740 2.400 2244.940 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1985.340 2.400 1986.540 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 571.620 2924.800 572.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.940 2.400 1728.140 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1468.540 2.400 1469.740 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1210.140 2.400 1211.340 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 951.740 2.400 952.940 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 693.340 2.400 694.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 434.940 2.400 436.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 241.140 2.400 242.340 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 47.340 2.400 48.540 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 769.500 2924.800 770.700 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1165.260 2924.800 1166.460 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1363.140 2924.800 1364.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1626.980 2924.800 1628.180 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1890.820 2924.800 1892.020 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2154.660 2924.800 2155.860 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 109.900 2924.800 111.100 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2352.540 2924.800 2353.740 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2616.380 2924.800 2617.580 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2880.220 2924.800 2881.420 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3144.060 2924.800 3145.260 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3407.900 2924.800 3409.100 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 3517.600 2714.970 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 3517.600 2391.130 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.730 3517.600 2067.290 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.890 3517.600 1743.450 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 307.780 2924.800 308.980 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.210 3517.600 1095.770 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.370 3517.600 771.930 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.530 3517.600 448.090 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 3517.600 124.250 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3341.940 2.400 3343.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3083.540 2.400 3084.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2825.140 2.400 2826.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2566.740 2.400 2567.940 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2308.340 2.400 2309.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2049.940 2.400 2051.140 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 505.660 2924.800 506.860 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1533.140 2.400 1534.340 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1274.740 2.400 1275.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1016.340 2.400 1017.540 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 757.940 2.400 759.140 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 499.540 2.400 500.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 305.740 2.400 306.940 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 111.940 2.400 113.140 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 703.540 2924.800 704.740 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 901.420 2924.800 902.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1099.300 2924.800 1100.500 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1297.180 2924.800 1298.380 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1561.020 2924.800 1562.220 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2088.700 2924.800 2089.900 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.970 -4.800 684.530 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.970 -4.800 2340.530 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.530 -4.800 2357.090 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.090 -4.800 2373.650 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.650 -4.800 2390.210 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2406.210 -4.800 2406.770 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.330 -4.800 2439.890 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.890 -4.800 2456.450 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.450 -4.800 2473.010 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.010 -4.800 2489.570 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.570 -4.800 850.130 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.570 -4.800 2506.130 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.130 -4.800 2522.690 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.690 -4.800 2539.250 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.250 -4.800 2555.810 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.370 -4.800 2588.930 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.930 -4.800 2605.490 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.490 -4.800 2622.050 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.050 -4.800 2638.610 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.610 -4.800 2655.170 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.130 -4.800 866.690 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.170 -4.800 2671.730 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.730 -4.800 2688.290 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.290 -4.800 2704.850 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.850 -4.800 2721.410 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.410 -4.800 2737.970 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.970 -4.800 2754.530 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.530 -4.800 2771.090 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.090 -4.800 2787.650 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.250 -4.800 899.810 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.810 -4.800 916.370 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 -4.800 932.930 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.930 -4.800 949.490 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.490 -4.800 966.050 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.050 -4.800 982.610 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.610 -4.800 999.170 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.530 -4.800 701.090 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.170 -4.800 1015.730 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.730 -4.800 1032.290 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.290 -4.800 1048.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.850 -4.800 1065.410 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.410 -4.800 1081.970 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.970 -4.800 1098.530 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.090 -4.800 1131.650 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.650 -4.800 1148.210 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.210 -4.800 1164.770 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.090 -4.800 717.650 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.770 -4.800 1181.330 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.330 -4.800 1197.890 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.890 -4.800 1214.450 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.450 -4.800 1231.010 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.010 -4.800 1247.570 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.570 -4.800 1264.130 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.130 -4.800 1280.690 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.690 -4.800 1297.250 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.250 -4.800 1313.810 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.810 -4.800 1330.370 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.650 -4.800 734.210 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.930 -4.800 1363.490 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.490 -4.800 1380.050 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.050 -4.800 1396.610 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.610 -4.800 1413.170 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.170 -4.800 1429.730 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.730 -4.800 1446.290 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.290 -4.800 1462.850 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.850 -4.800 1479.410 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.210 -4.800 750.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.970 -4.800 1512.530 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.530 -4.800 1529.090 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.650 -4.800 1562.210 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.210 -4.800 1578.770 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.770 -4.800 1595.330 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.330 -4.800 1611.890 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.450 -4.800 1645.010 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.010 -4.800 1661.570 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.770 -4.800 767.330 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.570 -4.800 1678.130 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.130 -4.800 1694.690 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 -4.800 1744.370 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.370 -4.800 1760.930 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.930 -4.800 1777.490 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.050 -4.800 1810.610 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.610 -4.800 1827.170 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.330 -4.800 783.890 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.170 -4.800 1843.730 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.730 -4.800 1860.290 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.850 -4.800 1893.410 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.410 -4.800 1909.970 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.970 -4.800 1926.530 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.530 -4.800 1943.090 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.650 -4.800 1976.210 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.210 -4.800 1992.770 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.890 -4.800 800.450 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.770 -4.800 2009.330 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.330 -4.800 2025.890 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.450 -4.800 2059.010 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.010 -4.800 2075.570 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.570 -4.800 2092.130 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.130 -4.800 2108.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.250 -4.800 2141.810 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.810 -4.800 2158.370 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.450 -4.800 817.010 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.370 -4.800 2174.930 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.050 -4.800 2224.610 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.610 -4.800 2241.170 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.730 -4.800 2274.290 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.850 -4.800 2307.410 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.410 -4.800 2323.970 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.010 -4.800 833.570 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.490 -4.800 690.050 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.050 -4.800 2362.610 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.170 -4.800 2395.730 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.730 -4.800 2412.290 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.290 -4.800 2428.850 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.850 -4.800 2445.410 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.970 -4.800 2478.530 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.090 -4.800 855.650 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.090 -4.800 2511.650 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.650 -4.800 2528.210 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.770 -4.800 2561.330 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.330 -4.800 2577.890 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.890 -4.800 2594.450 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.450 -4.800 2611.010 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.570 -4.800 2644.130 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.130 -4.800 2660.690 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.650 -4.800 872.210 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.690 -4.800 2677.250 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.250 -4.800 2693.810 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.930 -4.800 2743.490 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.490 -4.800 2760.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.050 -4.800 2776.610 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.210 -4.800 888.770 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.770 -4.800 905.330 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.330 -4.800 921.890 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.890 -4.800 938.450 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.450 -4.800 955.010 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.010 -4.800 971.570 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.570 -4.800 988.130 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.130 -4.800 1004.690 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.690 -4.800 1021.250 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.810 -4.800 1054.370 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.370 -4.800 1070.930 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.930 -4.800 1087.490 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.490 -4.800 1104.050 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.050 -4.800 1120.610 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.610 -4.800 1137.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.170 -4.800 1153.730 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.730 -4.800 1170.290 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.610 -4.800 723.170 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.290 -4.800 1186.850 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.850 -4.800 1203.410 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.410 -4.800 1219.970 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.970 -4.800 1236.530 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.530 -4.800 1253.090 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.650 -4.800 1286.210 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.210 -4.800 1302.770 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.770 -4.800 1319.330 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.330 -4.800 1335.890 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.170 -4.800 739.730 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.890 -4.800 1352.450 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.450 -4.800 1369.010 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.010 -4.800 1385.570 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.570 -4.800 1402.130 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.690 -4.800 1435.250 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.250 -4.800 1451.810 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.810 -4.800 1468.370 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.370 -4.800 1484.930 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.930 -4.800 1501.490 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.730 -4.800 756.290 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.490 -4.800 1518.050 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.050 -4.800 1534.610 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.610 -4.800 1551.170 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.170 -4.800 1567.730 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.730 -4.800 1584.290 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.290 -4.800 1600.850 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.850 -4.800 1617.410 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.410 -4.800 1633.970 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.530 -4.800 1667.090 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.290 -4.800 772.850 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.090 -4.800 1683.650 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.650 -4.800 1700.210 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.210 -4.800 1716.770 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.770 -4.800 1733.330 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.330 -4.800 1749.890 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.890 -4.800 1766.450 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.450 -4.800 1783.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.010 -4.800 1799.570 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.570 -4.800 1816.130 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.130 -4.800 1832.690 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.690 -4.800 1849.250 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.250 -4.800 1865.810 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.370 -4.800 1898.930 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.930 -4.800 1915.490 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.490 -4.800 1932.050 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.050 -4.800 1948.610 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.610 -4.800 1965.170 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.170 -4.800 1981.730 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.730 -4.800 1998.290 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.290 -4.800 2014.850 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.850 -4.800 2031.410 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.410 -4.800 2047.970 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.970 -4.800 2064.530 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.530 -4.800 2081.090 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.090 -4.800 2097.650 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.210 -4.800 2130.770 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.770 -4.800 2147.330 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.330 -4.800 2163.890 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.970 -4.800 822.530 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.890 -4.800 2180.450 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.450 -4.800 2197.010 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.570 -4.800 2230.130 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.130 -4.800 2246.690 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.690 -4.800 2263.250 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.250 -4.800 2279.810 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.370 -4.800 2312.930 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.930 -4.800 2329.490 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.530 -4.800 839.090 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.010 -4.800 695.570 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.010 -4.800 2351.570 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.570 -4.800 2368.130 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.130 -4.800 2384.690 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.690 -4.800 2401.250 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.810 -4.800 2434.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.370 -4.800 2450.930 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.930 -4.800 2467.490 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.490 -4.800 2484.050 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.050 -4.800 2500.610 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.610 -4.800 861.170 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.610 -4.800 2517.170 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.170 -4.800 2533.730 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.730 -4.800 2550.290 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.290 -4.800 2566.850 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.850 -4.800 2583.410 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.410 -4.800 2599.970 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.970 -4.800 2616.530 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.530 -4.800 2633.090 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.650 -4.800 2666.210 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.210 -4.800 2682.770 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.770 -4.800 2699.330 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.330 -4.800 2715.890 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2731.890 -4.800 2732.450 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.450 -4.800 2749.010 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.010 -4.800 2765.570 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.570 -4.800 2782.130 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 -4.800 2798.690 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.730 -4.800 894.290 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.290 -4.800 910.850 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.850 -4.800 927.410 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.410 -4.800 943.970 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.530 -4.800 977.090 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.090 -4.800 993.650 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.650 -4.800 1010.210 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.570 -4.800 712.130 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.210 -4.800 1026.770 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.330 -4.800 1059.890 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.890 -4.800 1076.450 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.450 -4.800 1093.010 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.010 -4.800 1109.570 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.130 -4.800 1142.690 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.690 -4.800 1159.250 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.250 -4.800 1175.810 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.930 -4.800 1225.490 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.490 -4.800 1242.050 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.050 -4.800 1258.610 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.610 -4.800 1275.170 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.730 -4.800 1308.290 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.290 -4.800 1324.850 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.850 -4.800 1341.410 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.690 -4.800 745.250 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.410 -4.800 1357.970 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.530 -4.800 1391.090 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.090 -4.800 1407.650 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.210 -4.800 1440.770 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.330 -4.800 1473.890 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.890 -4.800 1490.450 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.450 -4.800 1507.010 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.250 -4.800 761.810 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.010 -4.800 1523.570 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.130 -4.800 1556.690 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.250 -4.800 1589.810 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.810 -4.800 1606.370 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.370 -4.800 1622.930 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.930 -4.800 1639.490 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.490 -4.800 1656.050 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.050 -4.800 1672.610 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.810 -4.800 778.370 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.610 -4.800 1689.170 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.170 -4.800 1705.730 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.730 -4.800 1722.290 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.290 -4.800 1738.850 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.850 -4.800 1755.410 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.410 -4.800 1771.970 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.970 -4.800 1788.530 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.090 -4.800 1821.650 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.650 -4.800 1838.210 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.210 -4.800 1854.770 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.770 -4.800 1871.330 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.330 -4.800 1887.890 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.890 -4.800 1904.450 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.450 -4.800 1921.010 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.010 -4.800 1937.570 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.570 -4.800 1954.130 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.130 -4.800 1970.690 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.250 -4.800 2003.810 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.930 -4.800 811.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.810 -4.800 2020.370 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.930 -4.800 2053.490 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.490 -4.800 2070.050 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.050 -4.800 2086.610 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.610 -4.800 2103.170 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.170 -4.800 2119.730 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.730 -4.800 2136.290 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.290 -4.800 2152.850 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.850 -4.800 2169.410 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.490 -4.800 828.050 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.410 -4.800 2185.970 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.970 -4.800 2202.530 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.530 -4.800 2219.090 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.090 -4.800 2235.650 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.650 -4.800 2252.210 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.770 -4.800 2285.330 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.330 -4.800 2301.890 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.890 -4.800 2318.450 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.450 -4.800 2335.010 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.050 -4.800 844.610 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.170 -4.800 2809.730 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.690 -4.800 2815.250 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2820.210 -4.800 2820.770 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.970 -39.820 27.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.970 -39.820 127.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.970 1726.300 127.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.970 3440.300 127.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.970 -39.820 227.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.970 1726.300 227.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.970 3440.300 227.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 -39.820 327.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 1726.300 327.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 3440.300 327.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.970 -39.820 427.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.970 1726.300 427.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.970 3440.300 427.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.970 -39.820 527.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.970 1726.300 527.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.970 3440.300 527.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.970 -39.820 627.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.970 1726.300 627.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.970 3440.300 627.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.970 -39.820 727.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.970 1726.300 727.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.970 3440.300 727.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.970 -39.820 827.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.970 1726.300 827.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.970 3440.300 827.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.970 -39.820 927.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.970 1726.300 927.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.970 3440.300 927.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.970 -39.820 1027.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.970 1726.300 1027.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.970 3440.300 1027.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.970 -39.820 1127.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.970 1726.300 1127.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.970 3440.300 1127.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 -39.820 1227.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 1726.300 1227.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 3440.300 1227.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.970 -39.820 1327.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.970 1726.300 1327.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.970 3440.300 1327.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.970 -39.820 1427.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.970 -39.820 1527.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.970 1726.300 1527.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.970 3440.300 1527.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.970 -39.820 1627.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.970 1726.300 1627.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.970 3440.300 1627.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.970 -39.820 1727.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.970 1726.300 1727.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.970 3440.300 1727.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.970 -39.820 1827.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.970 1726.300 1827.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.970 3440.300 1827.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.970 -39.820 1927.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.970 1726.300 1927.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.970 3440.300 1927.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.970 -39.820 2027.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.970 1726.300 2027.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.970 3440.300 2027.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 -39.820 2127.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 1726.300 2127.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 3440.300 2127.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.970 -39.820 2227.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.970 1726.300 2227.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.970 3440.300 2227.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.970 -39.820 2327.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.970 1726.300 2327.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.970 3440.300 2327.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.970 -39.820 2427.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.970 1726.300 2427.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.970 3440.300 2427.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.970 -39.820 2527.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.970 1726.300 2527.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.970 3440.300 2527.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.970 -39.820 2627.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.970 1726.300 2627.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.970 3440.300 2627.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.970 -39.820 2727.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.970 1726.300 2727.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.970 3440.300 2727.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.970 -39.820 2827.070 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.970 1726.300 2827.070 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.970 3440.300 2827.070 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 29.330 2964.800 32.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 129.330 2964.800 132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 229.330 2964.800 232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 329.330 2964.800 332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 429.330 2964.800 432.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 529.330 2964.800 532.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 629.330 2964.800 632.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 729.330 2964.800 732.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 829.330 2964.800 832.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 929.330 2964.800 932.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1029.330 2964.800 1032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1129.330 2964.800 1132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1229.330 2964.800 1232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1329.330 2964.800 1332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1429.330 2964.800 1432.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1529.330 2964.800 1532.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1629.330 2964.800 1632.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1729.330 2964.800 1732.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1829.330 2964.800 1832.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1929.330 2964.800 1932.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2029.330 2964.800 2032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2129.330 2964.800 2132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2229.330 2964.800 2232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2329.330 2964.800 2332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2429.330 2964.800 2432.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2529.330 2964.800 2532.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2629.330 2964.800 2632.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2729.330 2964.800 2732.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2829.330 2964.800 2832.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2929.330 2964.800 2932.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3029.330 2964.800 3032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3129.330 2964.800 3132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3229.330 2964.800 3232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3329.330 2964.800 3332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3429.330 2964.800 3432.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2873.910 1814.000 2877.010 1825.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2873.910 100.400 2877.010 1730.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 2873.910 1825.760 2877.010 3443.760 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -21.180 -15.820 -18.080 3535.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 -15.820 2940.800 -12.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 3532.400 2940.800 3535.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2937.700 -15.820 2940.800 3535.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.170 -39.820 43.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.170 -39.820 143.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.170 3440.300 143.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 240.170 -39.820 243.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 240.170 3440.300 243.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 340.170 -39.820 343.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 340.170 3440.300 343.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 440.170 -39.820 443.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 440.170 3440.300 443.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 540.170 -39.820 543.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 540.170 3440.300 543.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 640.170 -39.820 643.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 640.170 3440.300 643.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 740.170 -39.820 743.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 740.170 3440.300 743.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.170 -39.820 843.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.170 3440.300 843.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 940.170 -39.820 943.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 940.170 3440.300 943.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1040.170 -39.820 1043.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1040.170 3440.300 1043.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1140.170 -39.820 1143.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1140.170 3440.300 1143.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1240.170 -39.820 1243.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1240.170 3440.300 1243.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.170 -39.820 1343.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.170 3440.300 1343.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1440.170 -39.820 1443.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1540.170 -39.820 1543.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1540.170 3440.300 1543.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.170 -39.820 1643.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.170 3440.300 1643.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1740.170 -39.820 1743.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1740.170 3440.300 1743.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1840.170 -39.820 1843.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1840.170 3440.300 1843.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1940.170 -39.820 1943.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1940.170 3440.300 1943.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2040.170 -39.820 2043.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2040.170 3440.300 2043.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2140.170 -39.820 2143.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2140.170 3440.300 2143.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.170 -39.820 2243.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.170 3440.300 2243.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2340.170 -39.820 2343.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2340.170 3440.300 2343.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2440.170 -39.820 2443.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2440.170 3440.300 2443.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2540.170 -39.820 2543.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2540.170 3440.300 2543.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2640.170 -39.820 2643.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2640.170 3440.300 2643.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2740.170 -39.820 2743.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2740.170 3440.300 2743.270 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.170 -39.820 2843.270 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.170 3440.300 2843.270 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 45.530 2964.800 48.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 145.530 2964.800 148.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 245.530 2964.800 248.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 345.530 2964.800 348.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 445.530 2964.800 448.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 545.530 2964.800 548.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 645.530 2964.800 648.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 745.530 2964.800 748.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 845.530 2964.800 848.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 945.530 2964.800 948.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1045.530 2964.800 1048.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1145.530 2964.800 1148.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1245.530 2964.800 1248.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1345.530 2964.800 1348.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1445.530 2964.800 1448.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1545.530 2964.800 1548.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1645.530 2964.800 1648.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1745.530 2964.800 1748.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1845.530 2964.800 1848.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1945.530 2964.800 1948.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2045.530 2964.800 2048.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2145.530 2964.800 2148.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2245.530 2964.800 2248.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2345.530 2964.800 2348.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2445.530 2964.800 2448.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2545.530 2964.800 2548.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2645.530 2964.800 2648.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2745.530 2964.800 2748.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2845.530 2964.800 2848.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2945.530 2964.800 2948.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3045.530 2964.800 3048.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3145.530 2964.800 3148.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3245.530 2964.800 3248.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3345.530 2964.800 3348.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3445.530 2964.800 3448.630 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -30.780 -25.420 -27.680 3545.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 -25.420 2950.400 -22.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 3542.000 2950.400 3545.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2947.300 -25.420 2950.400 3545.100 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -40.380 -35.020 -37.280 3554.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 -35.020 2960.000 -31.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 3551.600 2960.000 3554.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2956.900 -35.020 2960.000 3554.700 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -35.580 -30.220 -32.480 3549.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 -30.220 2955.200 -27.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 3546.800 2955.200 3549.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2952.100 -30.220 2955.200 3549.900 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -45.180 -39.820 -42.080 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 -39.820 2964.800 -36.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3556.400 2964.800 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2961.700 -39.820 2964.800 3559.500 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.070 -39.820 35.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.070 -39.820 135.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.070 1726.300 135.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.070 3440.300 135.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.070 -39.820 235.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.070 1726.300 235.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.070 3440.300 235.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.070 -39.820 335.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.070 1726.300 335.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.070 3440.300 335.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.070 -39.820 435.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.070 1726.300 435.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.070 3440.300 435.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.070 -39.820 535.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.070 1726.300 535.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.070 3440.300 535.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.070 -39.820 635.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.070 1726.300 635.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.070 3440.300 635.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.070 -39.820 735.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.070 1726.300 735.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.070 3440.300 735.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.070 -39.820 835.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.070 1726.300 835.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.070 3440.300 835.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.070 -39.820 935.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.070 1726.300 935.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.070 3440.300 935.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.070 -39.820 1035.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.070 1726.300 1035.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.070 3440.300 1035.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.070 -39.820 1135.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.070 1726.300 1135.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.070 3440.300 1135.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.070 -39.820 1235.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.070 1726.300 1235.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.070 3440.300 1235.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1332.070 -39.820 1335.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1332.070 1726.300 1335.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1332.070 3440.300 1335.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1432.070 -39.820 1435.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1532.070 -39.820 1535.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1532.070 1726.300 1535.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1532.070 3440.300 1535.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.070 -39.820 1635.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.070 1726.300 1635.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.070 3440.300 1635.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1732.070 -39.820 1735.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1732.070 1726.300 1735.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1732.070 3440.300 1735.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1832.070 -39.820 1835.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1832.070 1726.300 1835.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1832.070 3440.300 1835.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.070 -39.820 1935.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.070 1726.300 1935.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.070 3440.300 1935.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.070 -39.820 2035.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.070 1726.300 2035.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.070 3440.300 2035.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.070 -39.820 2135.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.070 1726.300 2135.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.070 3440.300 2135.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.070 -39.820 2235.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.070 1726.300 2235.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.070 3440.300 2235.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.070 -39.820 2335.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.070 1726.300 2335.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.070 3440.300 2335.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.070 -39.820 2435.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.070 1726.300 2435.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.070 3440.300 2435.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.070 -39.820 2535.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.070 1726.300 2535.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.070 3440.300 2535.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.070 -39.820 2635.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.070 1726.300 2635.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.070 3440.300 2635.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.070 -39.820 2735.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.070 1726.300 2735.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.070 3440.300 2735.170 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.070 -39.820 2835.170 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.070 1726.300 2835.170 1819.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.070 3440.300 2835.170 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 37.430 2964.800 40.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 137.430 2964.800 140.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 237.430 2964.800 240.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 337.430 2964.800 340.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 437.430 2964.800 440.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 537.430 2964.800 540.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 637.430 2964.800 640.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 737.430 2964.800 740.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 837.430 2964.800 840.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 937.430 2964.800 940.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1037.430 2964.800 1040.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1137.430 2964.800 1140.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1237.430 2964.800 1240.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1337.430 2964.800 1340.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1437.430 2964.800 1440.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1537.430 2964.800 1540.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1637.430 2964.800 1640.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1737.430 2964.800 1740.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1837.430 2964.800 1840.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1937.430 2964.800 1940.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2037.430 2964.800 2040.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2137.430 2964.800 2140.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2237.430 2964.800 2240.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2337.430 2964.800 2340.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2437.430 2964.800 2440.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2537.430 2964.800 2540.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2637.430 2964.800 2640.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2737.430 2964.800 2740.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2837.430 2964.800 2840.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2937.430 2964.800 2940.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3037.430 2964.800 3040.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3137.430 2964.800 3140.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3237.430 2964.800 3240.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3337.430 2964.800 3340.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3437.430 2964.800 3440.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 2882.190 1814.000 2885.290 1825.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2882.190 100.400 2885.290 1730.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 2882.190 1825.760 2885.290 3443.760 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -25.980 -20.620 -22.880 3540.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 -20.620 2945.600 -17.520 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 3537.200 2945.600 3540.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2942.500 -20.620 2945.600 3540.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.270 -39.820 51.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.270 -39.820 151.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.270 3440.300 151.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.270 -39.820 251.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.270 3440.300 251.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 348.270 -39.820 351.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 348.270 3440.300 351.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.270 -39.820 451.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.270 3440.300 451.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.270 -39.820 551.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.270 3440.300 551.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.270 -39.820 651.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.270 3440.300 651.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 748.270 -39.820 751.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 748.270 3440.300 751.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.270 -39.820 851.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.270 3440.300 851.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 948.270 -39.820 951.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 948.270 3440.300 951.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1048.270 -39.820 1051.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1048.270 3440.300 1051.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1148.270 -39.820 1151.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1148.270 3440.300 1151.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.270 -39.820 1251.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.270 3440.300 1251.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1348.270 -39.820 1351.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1348.270 3440.300 1351.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.270 -39.820 1451.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.270 -39.820 1551.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.270 3440.300 1551.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.270 -39.820 1651.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.270 3440.300 1651.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1748.270 -39.820 1751.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1748.270 3440.300 1751.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.270 -39.820 1851.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.270 3440.300 1851.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1948.270 -39.820 1951.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1948.270 3440.300 1951.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.270 -39.820 2051.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.270 3440.300 2051.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2148.270 -39.820 2151.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2148.270 3440.300 2151.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.270 -39.820 2251.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.270 3440.300 2251.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.270 -39.820 2351.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.270 3440.300 2351.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2448.270 -39.820 2451.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2448.270 3440.300 2451.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2548.270 -39.820 2551.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2548.270 3440.300 2551.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2648.270 -39.820 2651.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2648.270 3440.300 2651.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2748.270 -39.820 2751.370 105.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2748.270 3440.300 2751.370 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2848.270 -39.820 2851.370 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 53.630 2964.800 56.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 153.630 2964.800 156.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 253.630 2964.800 256.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 353.630 2964.800 356.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 453.630 2964.800 456.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 553.630 2964.800 556.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 653.630 2964.800 656.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 753.630 2964.800 756.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 853.630 2964.800 856.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 953.630 2964.800 956.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1053.630 2964.800 1056.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1153.630 2964.800 1156.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1253.630 2964.800 1256.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1353.630 2964.800 1356.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1453.630 2964.800 1456.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1553.630 2964.800 1556.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1653.630 2964.800 1656.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1753.630 2964.800 1756.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1853.630 2964.800 1856.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1953.630 2964.800 1956.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2053.630 2964.800 2056.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2153.630 2964.800 2156.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2253.630 2964.800 2256.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2353.630 2964.800 2356.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2453.630 2964.800 2456.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2553.630 2964.800 2556.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2653.630 2964.800 2656.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2753.630 2964.800 2756.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2853.630 2964.800 2856.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2953.630 2964.800 2956.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3053.630 2964.800 3056.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3153.630 2964.800 3156.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3253.630 2964.800 3256.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3353.630 2964.800 3356.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3453.630 2964.800 3456.730 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 -4.800 99.410 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 -4.800 104.930 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 -4.800 110.450 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 -4.800 320.210 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.210 -4.800 336.770 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.770 -4.800 353.330 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.330 -4.800 369.890 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.890 -4.800 386.450 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.450 -4.800 403.010 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.570 -4.800 436.130 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.130 -4.800 452.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.690 -4.800 469.250 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.050 -4.800 154.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.250 -4.800 485.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.810 -4.800 502.370 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.370 -4.800 518.930 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.930 -4.800 535.490 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.490 -4.800 552.050 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.050 -4.800 568.610 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.610 -4.800 585.170 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.170 -4.800 601.730 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.730 -4.800 618.290 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.290 -4.800 634.850 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.130 -4.800 176.690 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.410 -4.800 667.970 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.210 -4.800 198.770 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.290 -4.800 220.850 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.850 -4.800 237.410 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.410 -4.800 253.970 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 -4.800 287.090 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.090 -4.800 303.650 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.490 -4.800 138.050 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.170 -4.800 325.730 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.730 -4.800 342.290 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.290 -4.800 358.850 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.410 -4.800 391.970 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.970 -4.800 408.530 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.090 -4.800 441.650 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.210 -4.800 474.770 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.570 -4.800 160.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.770 -4.800 491.330 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.330 -4.800 507.890 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.890 -4.800 524.450 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.010 -4.800 557.570 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.130 -4.800 590.690 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.690 -4.800 607.250 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.810 -4.800 640.370 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.650 -4.800 182.210 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.370 -4.800 656.930 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.930 -4.800 673.490 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 -4.800 204.290 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.810 -4.800 226.370 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 -4.800 242.930 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.930 -4.800 259.490 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.490 -4.800 276.050 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.610 -4.800 309.170 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.010 -4.800 143.570 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.690 -4.800 331.250 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 -4.800 364.370 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.370 -4.800 380.930 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.930 -4.800 397.490 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.490 -4.800 414.050 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.050 -4.800 430.610 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.610 -4.800 447.170 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.170 -4.800 463.730 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.730 -4.800 480.290 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.090 -4.800 165.650 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.850 -4.800 513.410 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.410 -4.800 529.970 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.970 -4.800 546.530 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.530 -4.800 563.090 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.090 -4.800 579.650 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.650 -4.800 596.210 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.210 -4.800 612.770 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.770 -4.800 629.330 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.330 -4.800 645.890 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 -4.800 187.730 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.890 -4.800 662.450 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.450 -4.800 679.010 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 -4.800 231.890 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.890 -4.800 248.450 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 -4.800 265.010 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.010 -4.800 281.570 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 -4.800 298.130 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.130 -4.800 314.690 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530 -4.800 149.090 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.770 -4.800 215.330 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 5.520 4.120 2914.100 3509.040 ;
      LAYER met2 ;
        RECT 12.060 3517.320 42.450 3517.600 ;
        RECT 43.570 3517.320 123.410 3517.600 ;
        RECT 124.530 3517.320 204.370 3517.600 ;
        RECT 205.490 3517.320 285.330 3517.600 ;
        RECT 286.450 3517.320 366.290 3517.600 ;
        RECT 367.410 3517.320 447.250 3517.600 ;
        RECT 448.370 3517.320 528.210 3517.600 ;
        RECT 529.330 3517.320 609.170 3517.600 ;
        RECT 610.290 3517.320 690.130 3517.600 ;
        RECT 691.250 3517.320 771.090 3517.600 ;
        RECT 772.210 3517.320 852.050 3517.600 ;
        RECT 853.170 3517.320 933.010 3517.600 ;
        RECT 934.130 3517.320 1013.970 3517.600 ;
        RECT 1015.090 3517.320 1094.930 3517.600 ;
        RECT 1096.050 3517.320 1175.890 3517.600 ;
        RECT 1177.010 3517.320 1256.850 3517.600 ;
        RECT 1257.970 3517.320 1337.810 3517.600 ;
        RECT 1338.930 3517.320 1418.770 3517.600 ;
        RECT 1419.890 3517.320 1499.730 3517.600 ;
        RECT 1500.850 3517.320 1580.690 3517.600 ;
        RECT 1581.810 3517.320 1661.650 3517.600 ;
        RECT 1662.770 3517.320 1742.610 3517.600 ;
        RECT 1743.730 3517.320 1823.570 3517.600 ;
        RECT 1824.690 3517.320 1904.530 3517.600 ;
        RECT 1905.650 3517.320 1985.490 3517.600 ;
        RECT 1986.610 3517.320 2066.450 3517.600 ;
        RECT 2067.570 3517.320 2147.410 3517.600 ;
        RECT 2148.530 3517.320 2228.370 3517.600 ;
        RECT 2229.490 3517.320 2309.330 3517.600 ;
        RECT 2310.450 3517.320 2390.290 3517.600 ;
        RECT 2391.410 3517.320 2471.250 3517.600 ;
        RECT 2472.370 3517.320 2552.210 3517.600 ;
        RECT 2553.330 3517.320 2633.170 3517.600 ;
        RECT 2634.290 3517.320 2714.130 3517.600 ;
        RECT 2715.250 3517.320 2795.090 3517.600 ;
        RECT 2796.210 3517.320 2876.050 3517.600 ;
        RECT 2877.170 3517.320 2908.490 3517.600 ;
        RECT 12.060 2.680 2908.490 3517.320 ;
        RECT 12.060 0.950 98.570 2.680 ;
        RECT 99.690 0.950 104.090 2.680 ;
        RECT 105.210 0.950 109.610 2.680 ;
        RECT 110.730 0.950 115.130 2.680 ;
        RECT 116.250 0.950 120.650 2.680 ;
        RECT 121.770 0.950 126.170 2.680 ;
        RECT 127.290 0.950 131.690 2.680 ;
        RECT 132.810 0.950 137.210 2.680 ;
        RECT 138.330 0.950 142.730 2.680 ;
        RECT 143.850 0.950 148.250 2.680 ;
        RECT 149.370 0.950 153.770 2.680 ;
        RECT 154.890 0.950 159.290 2.680 ;
        RECT 160.410 0.950 164.810 2.680 ;
        RECT 165.930 0.950 170.330 2.680 ;
        RECT 171.450 0.950 175.850 2.680 ;
        RECT 176.970 0.950 181.370 2.680 ;
        RECT 182.490 0.950 186.890 2.680 ;
        RECT 188.010 0.950 192.410 2.680 ;
        RECT 193.530 0.950 197.930 2.680 ;
        RECT 199.050 0.950 203.450 2.680 ;
        RECT 204.570 0.950 208.970 2.680 ;
        RECT 210.090 0.950 214.490 2.680 ;
        RECT 215.610 0.950 220.010 2.680 ;
        RECT 221.130 0.950 225.530 2.680 ;
        RECT 226.650 0.950 231.050 2.680 ;
        RECT 232.170 0.950 236.570 2.680 ;
        RECT 237.690 0.950 242.090 2.680 ;
        RECT 243.210 0.950 247.610 2.680 ;
        RECT 248.730 0.950 253.130 2.680 ;
        RECT 254.250 0.950 258.650 2.680 ;
        RECT 259.770 0.950 264.170 2.680 ;
        RECT 265.290 0.950 269.690 2.680 ;
        RECT 270.810 0.950 275.210 2.680 ;
        RECT 276.330 0.950 280.730 2.680 ;
        RECT 281.850 0.950 286.250 2.680 ;
        RECT 287.370 0.950 291.770 2.680 ;
        RECT 292.890 0.950 297.290 2.680 ;
        RECT 298.410 0.950 302.810 2.680 ;
        RECT 303.930 0.950 308.330 2.680 ;
        RECT 309.450 0.950 313.850 2.680 ;
        RECT 314.970 0.950 319.370 2.680 ;
        RECT 320.490 0.950 324.890 2.680 ;
        RECT 326.010 0.950 330.410 2.680 ;
        RECT 331.530 0.950 335.930 2.680 ;
        RECT 337.050 0.950 341.450 2.680 ;
        RECT 342.570 0.950 346.970 2.680 ;
        RECT 348.090 0.950 352.490 2.680 ;
        RECT 353.610 0.950 358.010 2.680 ;
        RECT 359.130 0.950 363.530 2.680 ;
        RECT 364.650 0.950 369.050 2.680 ;
        RECT 370.170 0.950 374.570 2.680 ;
        RECT 375.690 0.950 380.090 2.680 ;
        RECT 381.210 0.950 385.610 2.680 ;
        RECT 386.730 0.950 391.130 2.680 ;
        RECT 392.250 0.950 396.650 2.680 ;
        RECT 397.770 0.950 402.170 2.680 ;
        RECT 403.290 0.950 407.690 2.680 ;
        RECT 408.810 0.950 413.210 2.680 ;
        RECT 414.330 0.950 418.730 2.680 ;
        RECT 419.850 0.950 424.250 2.680 ;
        RECT 425.370 0.950 429.770 2.680 ;
        RECT 430.890 0.950 435.290 2.680 ;
        RECT 436.410 0.950 440.810 2.680 ;
        RECT 441.930 0.950 446.330 2.680 ;
        RECT 447.450 0.950 451.850 2.680 ;
        RECT 452.970 0.950 457.370 2.680 ;
        RECT 458.490 0.950 462.890 2.680 ;
        RECT 464.010 0.950 468.410 2.680 ;
        RECT 469.530 0.950 473.930 2.680 ;
        RECT 475.050 0.950 479.450 2.680 ;
        RECT 480.570 0.950 484.970 2.680 ;
        RECT 486.090 0.950 490.490 2.680 ;
        RECT 491.610 0.950 496.010 2.680 ;
        RECT 497.130 0.950 501.530 2.680 ;
        RECT 502.650 0.950 507.050 2.680 ;
        RECT 508.170 0.950 512.570 2.680 ;
        RECT 513.690 0.950 518.090 2.680 ;
        RECT 519.210 0.950 523.610 2.680 ;
        RECT 524.730 0.950 529.130 2.680 ;
        RECT 530.250 0.950 534.650 2.680 ;
        RECT 535.770 0.950 540.170 2.680 ;
        RECT 541.290 0.950 545.690 2.680 ;
        RECT 546.810 0.950 551.210 2.680 ;
        RECT 552.330 0.950 556.730 2.680 ;
        RECT 557.850 0.950 562.250 2.680 ;
        RECT 563.370 0.950 567.770 2.680 ;
        RECT 568.890 0.950 573.290 2.680 ;
        RECT 574.410 0.950 578.810 2.680 ;
        RECT 579.930 0.950 584.330 2.680 ;
        RECT 585.450 0.950 589.850 2.680 ;
        RECT 590.970 0.950 595.370 2.680 ;
        RECT 596.490 0.950 600.890 2.680 ;
        RECT 602.010 0.950 606.410 2.680 ;
        RECT 607.530 0.950 611.930 2.680 ;
        RECT 613.050 0.950 617.450 2.680 ;
        RECT 618.570 0.950 622.970 2.680 ;
        RECT 624.090 0.950 628.490 2.680 ;
        RECT 629.610 0.950 634.010 2.680 ;
        RECT 635.130 0.950 639.530 2.680 ;
        RECT 640.650 0.950 645.050 2.680 ;
        RECT 646.170 0.950 650.570 2.680 ;
        RECT 651.690 0.950 656.090 2.680 ;
        RECT 657.210 0.950 661.610 2.680 ;
        RECT 662.730 0.950 667.130 2.680 ;
        RECT 668.250 0.950 672.650 2.680 ;
        RECT 673.770 0.950 678.170 2.680 ;
        RECT 679.290 0.950 683.690 2.680 ;
        RECT 684.810 0.950 689.210 2.680 ;
        RECT 690.330 0.950 694.730 2.680 ;
        RECT 695.850 0.950 700.250 2.680 ;
        RECT 701.370 0.950 705.770 2.680 ;
        RECT 706.890 0.950 711.290 2.680 ;
        RECT 712.410 0.950 716.810 2.680 ;
        RECT 717.930 0.950 722.330 2.680 ;
        RECT 723.450 0.950 727.850 2.680 ;
        RECT 728.970 0.950 733.370 2.680 ;
        RECT 734.490 0.950 738.890 2.680 ;
        RECT 740.010 0.950 744.410 2.680 ;
        RECT 745.530 0.950 749.930 2.680 ;
        RECT 751.050 0.950 755.450 2.680 ;
        RECT 756.570 0.950 760.970 2.680 ;
        RECT 762.090 0.950 766.490 2.680 ;
        RECT 767.610 0.950 772.010 2.680 ;
        RECT 773.130 0.950 777.530 2.680 ;
        RECT 778.650 0.950 783.050 2.680 ;
        RECT 784.170 0.950 788.570 2.680 ;
        RECT 789.690 0.950 794.090 2.680 ;
        RECT 795.210 0.950 799.610 2.680 ;
        RECT 800.730 0.950 805.130 2.680 ;
        RECT 806.250 0.950 810.650 2.680 ;
        RECT 811.770 0.950 816.170 2.680 ;
        RECT 817.290 0.950 821.690 2.680 ;
        RECT 822.810 0.950 827.210 2.680 ;
        RECT 828.330 0.950 832.730 2.680 ;
        RECT 833.850 0.950 838.250 2.680 ;
        RECT 839.370 0.950 843.770 2.680 ;
        RECT 844.890 0.950 849.290 2.680 ;
        RECT 850.410 0.950 854.810 2.680 ;
        RECT 855.930 0.950 860.330 2.680 ;
        RECT 861.450 0.950 865.850 2.680 ;
        RECT 866.970 0.950 871.370 2.680 ;
        RECT 872.490 0.950 876.890 2.680 ;
        RECT 878.010 0.950 882.410 2.680 ;
        RECT 883.530 0.950 887.930 2.680 ;
        RECT 889.050 0.950 893.450 2.680 ;
        RECT 894.570 0.950 898.970 2.680 ;
        RECT 900.090 0.950 904.490 2.680 ;
        RECT 905.610 0.950 910.010 2.680 ;
        RECT 911.130 0.950 915.530 2.680 ;
        RECT 916.650 0.950 921.050 2.680 ;
        RECT 922.170 0.950 926.570 2.680 ;
        RECT 927.690 0.950 932.090 2.680 ;
        RECT 933.210 0.950 937.610 2.680 ;
        RECT 938.730 0.950 943.130 2.680 ;
        RECT 944.250 0.950 948.650 2.680 ;
        RECT 949.770 0.950 954.170 2.680 ;
        RECT 955.290 0.950 959.690 2.680 ;
        RECT 960.810 0.950 965.210 2.680 ;
        RECT 966.330 0.950 970.730 2.680 ;
        RECT 971.850 0.950 976.250 2.680 ;
        RECT 977.370 0.950 981.770 2.680 ;
        RECT 982.890 0.950 987.290 2.680 ;
        RECT 988.410 0.950 992.810 2.680 ;
        RECT 993.930 0.950 998.330 2.680 ;
        RECT 999.450 0.950 1003.850 2.680 ;
        RECT 1004.970 0.950 1009.370 2.680 ;
        RECT 1010.490 0.950 1014.890 2.680 ;
        RECT 1016.010 0.950 1020.410 2.680 ;
        RECT 1021.530 0.950 1025.930 2.680 ;
        RECT 1027.050 0.950 1031.450 2.680 ;
        RECT 1032.570 0.950 1036.970 2.680 ;
        RECT 1038.090 0.950 1042.490 2.680 ;
        RECT 1043.610 0.950 1048.010 2.680 ;
        RECT 1049.130 0.950 1053.530 2.680 ;
        RECT 1054.650 0.950 1059.050 2.680 ;
        RECT 1060.170 0.950 1064.570 2.680 ;
        RECT 1065.690 0.950 1070.090 2.680 ;
        RECT 1071.210 0.950 1075.610 2.680 ;
        RECT 1076.730 0.950 1081.130 2.680 ;
        RECT 1082.250 0.950 1086.650 2.680 ;
        RECT 1087.770 0.950 1092.170 2.680 ;
        RECT 1093.290 0.950 1097.690 2.680 ;
        RECT 1098.810 0.950 1103.210 2.680 ;
        RECT 1104.330 0.950 1108.730 2.680 ;
        RECT 1109.850 0.950 1114.250 2.680 ;
        RECT 1115.370 0.950 1119.770 2.680 ;
        RECT 1120.890 0.950 1125.290 2.680 ;
        RECT 1126.410 0.950 1130.810 2.680 ;
        RECT 1131.930 0.950 1136.330 2.680 ;
        RECT 1137.450 0.950 1141.850 2.680 ;
        RECT 1142.970 0.950 1147.370 2.680 ;
        RECT 1148.490 0.950 1152.890 2.680 ;
        RECT 1154.010 0.950 1158.410 2.680 ;
        RECT 1159.530 0.950 1163.930 2.680 ;
        RECT 1165.050 0.950 1169.450 2.680 ;
        RECT 1170.570 0.950 1174.970 2.680 ;
        RECT 1176.090 0.950 1180.490 2.680 ;
        RECT 1181.610 0.950 1186.010 2.680 ;
        RECT 1187.130 0.950 1191.530 2.680 ;
        RECT 1192.650 0.950 1197.050 2.680 ;
        RECT 1198.170 0.950 1202.570 2.680 ;
        RECT 1203.690 0.950 1208.090 2.680 ;
        RECT 1209.210 0.950 1213.610 2.680 ;
        RECT 1214.730 0.950 1219.130 2.680 ;
        RECT 1220.250 0.950 1224.650 2.680 ;
        RECT 1225.770 0.950 1230.170 2.680 ;
        RECT 1231.290 0.950 1235.690 2.680 ;
        RECT 1236.810 0.950 1241.210 2.680 ;
        RECT 1242.330 0.950 1246.730 2.680 ;
        RECT 1247.850 0.950 1252.250 2.680 ;
        RECT 1253.370 0.950 1257.770 2.680 ;
        RECT 1258.890 0.950 1263.290 2.680 ;
        RECT 1264.410 0.950 1268.810 2.680 ;
        RECT 1269.930 0.950 1274.330 2.680 ;
        RECT 1275.450 0.950 1279.850 2.680 ;
        RECT 1280.970 0.950 1285.370 2.680 ;
        RECT 1286.490 0.950 1290.890 2.680 ;
        RECT 1292.010 0.950 1296.410 2.680 ;
        RECT 1297.530 0.950 1301.930 2.680 ;
        RECT 1303.050 0.950 1307.450 2.680 ;
        RECT 1308.570 0.950 1312.970 2.680 ;
        RECT 1314.090 0.950 1318.490 2.680 ;
        RECT 1319.610 0.950 1324.010 2.680 ;
        RECT 1325.130 0.950 1329.530 2.680 ;
        RECT 1330.650 0.950 1335.050 2.680 ;
        RECT 1336.170 0.950 1340.570 2.680 ;
        RECT 1341.690 0.950 1346.090 2.680 ;
        RECT 1347.210 0.950 1351.610 2.680 ;
        RECT 1352.730 0.950 1357.130 2.680 ;
        RECT 1358.250 0.950 1362.650 2.680 ;
        RECT 1363.770 0.950 1368.170 2.680 ;
        RECT 1369.290 0.950 1373.690 2.680 ;
        RECT 1374.810 0.950 1379.210 2.680 ;
        RECT 1380.330 0.950 1384.730 2.680 ;
        RECT 1385.850 0.950 1390.250 2.680 ;
        RECT 1391.370 0.950 1395.770 2.680 ;
        RECT 1396.890 0.950 1401.290 2.680 ;
        RECT 1402.410 0.950 1406.810 2.680 ;
        RECT 1407.930 0.950 1412.330 2.680 ;
        RECT 1413.450 0.950 1417.850 2.680 ;
        RECT 1418.970 0.950 1423.370 2.680 ;
        RECT 1424.490 0.950 1428.890 2.680 ;
        RECT 1430.010 0.950 1434.410 2.680 ;
        RECT 1435.530 0.950 1439.930 2.680 ;
        RECT 1441.050 0.950 1445.450 2.680 ;
        RECT 1446.570 0.950 1450.970 2.680 ;
        RECT 1452.090 0.950 1456.490 2.680 ;
        RECT 1457.610 0.950 1462.010 2.680 ;
        RECT 1463.130 0.950 1467.530 2.680 ;
        RECT 1468.650 0.950 1473.050 2.680 ;
        RECT 1474.170 0.950 1478.570 2.680 ;
        RECT 1479.690 0.950 1484.090 2.680 ;
        RECT 1485.210 0.950 1489.610 2.680 ;
        RECT 1490.730 0.950 1495.130 2.680 ;
        RECT 1496.250 0.950 1500.650 2.680 ;
        RECT 1501.770 0.950 1506.170 2.680 ;
        RECT 1507.290 0.950 1511.690 2.680 ;
        RECT 1512.810 0.950 1517.210 2.680 ;
        RECT 1518.330 0.950 1522.730 2.680 ;
        RECT 1523.850 0.950 1528.250 2.680 ;
        RECT 1529.370 0.950 1533.770 2.680 ;
        RECT 1534.890 0.950 1539.290 2.680 ;
        RECT 1540.410 0.950 1544.810 2.680 ;
        RECT 1545.930 0.950 1550.330 2.680 ;
        RECT 1551.450 0.950 1555.850 2.680 ;
        RECT 1556.970 0.950 1561.370 2.680 ;
        RECT 1562.490 0.950 1566.890 2.680 ;
        RECT 1568.010 0.950 1572.410 2.680 ;
        RECT 1573.530 0.950 1577.930 2.680 ;
        RECT 1579.050 0.950 1583.450 2.680 ;
        RECT 1584.570 0.950 1588.970 2.680 ;
        RECT 1590.090 0.950 1594.490 2.680 ;
        RECT 1595.610 0.950 1600.010 2.680 ;
        RECT 1601.130 0.950 1605.530 2.680 ;
        RECT 1606.650 0.950 1611.050 2.680 ;
        RECT 1612.170 0.950 1616.570 2.680 ;
        RECT 1617.690 0.950 1622.090 2.680 ;
        RECT 1623.210 0.950 1627.610 2.680 ;
        RECT 1628.730 0.950 1633.130 2.680 ;
        RECT 1634.250 0.950 1638.650 2.680 ;
        RECT 1639.770 0.950 1644.170 2.680 ;
        RECT 1645.290 0.950 1649.690 2.680 ;
        RECT 1650.810 0.950 1655.210 2.680 ;
        RECT 1656.330 0.950 1660.730 2.680 ;
        RECT 1661.850 0.950 1666.250 2.680 ;
        RECT 1667.370 0.950 1671.770 2.680 ;
        RECT 1672.890 0.950 1677.290 2.680 ;
        RECT 1678.410 0.950 1682.810 2.680 ;
        RECT 1683.930 0.950 1688.330 2.680 ;
        RECT 1689.450 0.950 1693.850 2.680 ;
        RECT 1694.970 0.950 1699.370 2.680 ;
        RECT 1700.490 0.950 1704.890 2.680 ;
        RECT 1706.010 0.950 1710.410 2.680 ;
        RECT 1711.530 0.950 1715.930 2.680 ;
        RECT 1717.050 0.950 1721.450 2.680 ;
        RECT 1722.570 0.950 1726.970 2.680 ;
        RECT 1728.090 0.950 1732.490 2.680 ;
        RECT 1733.610 0.950 1738.010 2.680 ;
        RECT 1739.130 0.950 1743.530 2.680 ;
        RECT 1744.650 0.950 1749.050 2.680 ;
        RECT 1750.170 0.950 1754.570 2.680 ;
        RECT 1755.690 0.950 1760.090 2.680 ;
        RECT 1761.210 0.950 1765.610 2.680 ;
        RECT 1766.730 0.950 1771.130 2.680 ;
        RECT 1772.250 0.950 1776.650 2.680 ;
        RECT 1777.770 0.950 1782.170 2.680 ;
        RECT 1783.290 0.950 1787.690 2.680 ;
        RECT 1788.810 0.950 1793.210 2.680 ;
        RECT 1794.330 0.950 1798.730 2.680 ;
        RECT 1799.850 0.950 1804.250 2.680 ;
        RECT 1805.370 0.950 1809.770 2.680 ;
        RECT 1810.890 0.950 1815.290 2.680 ;
        RECT 1816.410 0.950 1820.810 2.680 ;
        RECT 1821.930 0.950 1826.330 2.680 ;
        RECT 1827.450 0.950 1831.850 2.680 ;
        RECT 1832.970 0.950 1837.370 2.680 ;
        RECT 1838.490 0.950 1842.890 2.680 ;
        RECT 1844.010 0.950 1848.410 2.680 ;
        RECT 1849.530 0.950 1853.930 2.680 ;
        RECT 1855.050 0.950 1859.450 2.680 ;
        RECT 1860.570 0.950 1864.970 2.680 ;
        RECT 1866.090 0.950 1870.490 2.680 ;
        RECT 1871.610 0.950 1876.010 2.680 ;
        RECT 1877.130 0.950 1881.530 2.680 ;
        RECT 1882.650 0.950 1887.050 2.680 ;
        RECT 1888.170 0.950 1892.570 2.680 ;
        RECT 1893.690 0.950 1898.090 2.680 ;
        RECT 1899.210 0.950 1903.610 2.680 ;
        RECT 1904.730 0.950 1909.130 2.680 ;
        RECT 1910.250 0.950 1914.650 2.680 ;
        RECT 1915.770 0.950 1920.170 2.680 ;
        RECT 1921.290 0.950 1925.690 2.680 ;
        RECT 1926.810 0.950 1931.210 2.680 ;
        RECT 1932.330 0.950 1936.730 2.680 ;
        RECT 1937.850 0.950 1942.250 2.680 ;
        RECT 1943.370 0.950 1947.770 2.680 ;
        RECT 1948.890 0.950 1953.290 2.680 ;
        RECT 1954.410 0.950 1958.810 2.680 ;
        RECT 1959.930 0.950 1964.330 2.680 ;
        RECT 1965.450 0.950 1969.850 2.680 ;
        RECT 1970.970 0.950 1975.370 2.680 ;
        RECT 1976.490 0.950 1980.890 2.680 ;
        RECT 1982.010 0.950 1986.410 2.680 ;
        RECT 1987.530 0.950 1991.930 2.680 ;
        RECT 1993.050 0.950 1997.450 2.680 ;
        RECT 1998.570 0.950 2002.970 2.680 ;
        RECT 2004.090 0.950 2008.490 2.680 ;
        RECT 2009.610 0.950 2014.010 2.680 ;
        RECT 2015.130 0.950 2019.530 2.680 ;
        RECT 2020.650 0.950 2025.050 2.680 ;
        RECT 2026.170 0.950 2030.570 2.680 ;
        RECT 2031.690 0.950 2036.090 2.680 ;
        RECT 2037.210 0.950 2041.610 2.680 ;
        RECT 2042.730 0.950 2047.130 2.680 ;
        RECT 2048.250 0.950 2052.650 2.680 ;
        RECT 2053.770 0.950 2058.170 2.680 ;
        RECT 2059.290 0.950 2063.690 2.680 ;
        RECT 2064.810 0.950 2069.210 2.680 ;
        RECT 2070.330 0.950 2074.730 2.680 ;
        RECT 2075.850 0.950 2080.250 2.680 ;
        RECT 2081.370 0.950 2085.770 2.680 ;
        RECT 2086.890 0.950 2091.290 2.680 ;
        RECT 2092.410 0.950 2096.810 2.680 ;
        RECT 2097.930 0.950 2102.330 2.680 ;
        RECT 2103.450 0.950 2107.850 2.680 ;
        RECT 2108.970 0.950 2113.370 2.680 ;
        RECT 2114.490 0.950 2118.890 2.680 ;
        RECT 2120.010 0.950 2124.410 2.680 ;
        RECT 2125.530 0.950 2129.930 2.680 ;
        RECT 2131.050 0.950 2135.450 2.680 ;
        RECT 2136.570 0.950 2140.970 2.680 ;
        RECT 2142.090 0.950 2146.490 2.680 ;
        RECT 2147.610 0.950 2152.010 2.680 ;
        RECT 2153.130 0.950 2157.530 2.680 ;
        RECT 2158.650 0.950 2163.050 2.680 ;
        RECT 2164.170 0.950 2168.570 2.680 ;
        RECT 2169.690 0.950 2174.090 2.680 ;
        RECT 2175.210 0.950 2179.610 2.680 ;
        RECT 2180.730 0.950 2185.130 2.680 ;
        RECT 2186.250 0.950 2190.650 2.680 ;
        RECT 2191.770 0.950 2196.170 2.680 ;
        RECT 2197.290 0.950 2201.690 2.680 ;
        RECT 2202.810 0.950 2207.210 2.680 ;
        RECT 2208.330 0.950 2212.730 2.680 ;
        RECT 2213.850 0.950 2218.250 2.680 ;
        RECT 2219.370 0.950 2223.770 2.680 ;
        RECT 2224.890 0.950 2229.290 2.680 ;
        RECT 2230.410 0.950 2234.810 2.680 ;
        RECT 2235.930 0.950 2240.330 2.680 ;
        RECT 2241.450 0.950 2245.850 2.680 ;
        RECT 2246.970 0.950 2251.370 2.680 ;
        RECT 2252.490 0.950 2256.890 2.680 ;
        RECT 2258.010 0.950 2262.410 2.680 ;
        RECT 2263.530 0.950 2267.930 2.680 ;
        RECT 2269.050 0.950 2273.450 2.680 ;
        RECT 2274.570 0.950 2278.970 2.680 ;
        RECT 2280.090 0.950 2284.490 2.680 ;
        RECT 2285.610 0.950 2290.010 2.680 ;
        RECT 2291.130 0.950 2295.530 2.680 ;
        RECT 2296.650 0.950 2301.050 2.680 ;
        RECT 2302.170 0.950 2306.570 2.680 ;
        RECT 2307.690 0.950 2312.090 2.680 ;
        RECT 2313.210 0.950 2317.610 2.680 ;
        RECT 2318.730 0.950 2323.130 2.680 ;
        RECT 2324.250 0.950 2328.650 2.680 ;
        RECT 2329.770 0.950 2334.170 2.680 ;
        RECT 2335.290 0.950 2339.690 2.680 ;
        RECT 2340.810 0.950 2345.210 2.680 ;
        RECT 2346.330 0.950 2350.730 2.680 ;
        RECT 2351.850 0.950 2356.250 2.680 ;
        RECT 2357.370 0.950 2361.770 2.680 ;
        RECT 2362.890 0.950 2367.290 2.680 ;
        RECT 2368.410 0.950 2372.810 2.680 ;
        RECT 2373.930 0.950 2378.330 2.680 ;
        RECT 2379.450 0.950 2383.850 2.680 ;
        RECT 2384.970 0.950 2389.370 2.680 ;
        RECT 2390.490 0.950 2394.890 2.680 ;
        RECT 2396.010 0.950 2400.410 2.680 ;
        RECT 2401.530 0.950 2405.930 2.680 ;
        RECT 2407.050 0.950 2411.450 2.680 ;
        RECT 2412.570 0.950 2416.970 2.680 ;
        RECT 2418.090 0.950 2422.490 2.680 ;
        RECT 2423.610 0.950 2428.010 2.680 ;
        RECT 2429.130 0.950 2433.530 2.680 ;
        RECT 2434.650 0.950 2439.050 2.680 ;
        RECT 2440.170 0.950 2444.570 2.680 ;
        RECT 2445.690 0.950 2450.090 2.680 ;
        RECT 2451.210 0.950 2455.610 2.680 ;
        RECT 2456.730 0.950 2461.130 2.680 ;
        RECT 2462.250 0.950 2466.650 2.680 ;
        RECT 2467.770 0.950 2472.170 2.680 ;
        RECT 2473.290 0.950 2477.690 2.680 ;
        RECT 2478.810 0.950 2483.210 2.680 ;
        RECT 2484.330 0.950 2488.730 2.680 ;
        RECT 2489.850 0.950 2494.250 2.680 ;
        RECT 2495.370 0.950 2499.770 2.680 ;
        RECT 2500.890 0.950 2505.290 2.680 ;
        RECT 2506.410 0.950 2510.810 2.680 ;
        RECT 2511.930 0.950 2516.330 2.680 ;
        RECT 2517.450 0.950 2521.850 2.680 ;
        RECT 2522.970 0.950 2527.370 2.680 ;
        RECT 2528.490 0.950 2532.890 2.680 ;
        RECT 2534.010 0.950 2538.410 2.680 ;
        RECT 2539.530 0.950 2543.930 2.680 ;
        RECT 2545.050 0.950 2549.450 2.680 ;
        RECT 2550.570 0.950 2554.970 2.680 ;
        RECT 2556.090 0.950 2560.490 2.680 ;
        RECT 2561.610 0.950 2566.010 2.680 ;
        RECT 2567.130 0.950 2571.530 2.680 ;
        RECT 2572.650 0.950 2577.050 2.680 ;
        RECT 2578.170 0.950 2582.570 2.680 ;
        RECT 2583.690 0.950 2588.090 2.680 ;
        RECT 2589.210 0.950 2593.610 2.680 ;
        RECT 2594.730 0.950 2599.130 2.680 ;
        RECT 2600.250 0.950 2604.650 2.680 ;
        RECT 2605.770 0.950 2610.170 2.680 ;
        RECT 2611.290 0.950 2615.690 2.680 ;
        RECT 2616.810 0.950 2621.210 2.680 ;
        RECT 2622.330 0.950 2626.730 2.680 ;
        RECT 2627.850 0.950 2632.250 2.680 ;
        RECT 2633.370 0.950 2637.770 2.680 ;
        RECT 2638.890 0.950 2643.290 2.680 ;
        RECT 2644.410 0.950 2648.810 2.680 ;
        RECT 2649.930 0.950 2654.330 2.680 ;
        RECT 2655.450 0.950 2659.850 2.680 ;
        RECT 2660.970 0.950 2665.370 2.680 ;
        RECT 2666.490 0.950 2670.890 2.680 ;
        RECT 2672.010 0.950 2676.410 2.680 ;
        RECT 2677.530 0.950 2681.930 2.680 ;
        RECT 2683.050 0.950 2687.450 2.680 ;
        RECT 2688.570 0.950 2692.970 2.680 ;
        RECT 2694.090 0.950 2698.490 2.680 ;
        RECT 2699.610 0.950 2704.010 2.680 ;
        RECT 2705.130 0.950 2709.530 2.680 ;
        RECT 2710.650 0.950 2715.050 2.680 ;
        RECT 2716.170 0.950 2720.570 2.680 ;
        RECT 2721.690 0.950 2726.090 2.680 ;
        RECT 2727.210 0.950 2731.610 2.680 ;
        RECT 2732.730 0.950 2737.130 2.680 ;
        RECT 2738.250 0.950 2742.650 2.680 ;
        RECT 2743.770 0.950 2748.170 2.680 ;
        RECT 2749.290 0.950 2753.690 2.680 ;
        RECT 2754.810 0.950 2759.210 2.680 ;
        RECT 2760.330 0.950 2764.730 2.680 ;
        RECT 2765.850 0.950 2770.250 2.680 ;
        RECT 2771.370 0.950 2775.770 2.680 ;
        RECT 2776.890 0.950 2781.290 2.680 ;
        RECT 2782.410 0.950 2786.810 2.680 ;
        RECT 2787.930 0.950 2792.330 2.680 ;
        RECT 2793.450 0.950 2797.850 2.680 ;
        RECT 2798.970 0.950 2803.370 2.680 ;
        RECT 2804.490 0.950 2808.890 2.680 ;
        RECT 2810.010 0.950 2814.410 2.680 ;
        RECT 2815.530 0.950 2819.930 2.680 ;
        RECT 2821.050 0.950 2908.490 2.680 ;
      LAYER met3 ;
        RECT 2.400 3475.460 2917.600 3508.965 ;
        RECT 2.400 3473.460 2917.200 3475.460 ;
        RECT 2.400 3472.740 2917.600 3473.460 ;
        RECT 2.800 3470.740 2917.600 3472.740 ;
        RECT 2.400 3409.500 2917.600 3470.740 ;
        RECT 2.400 3408.140 2917.200 3409.500 ;
        RECT 2.800 3407.500 2917.200 3408.140 ;
        RECT 2.800 3406.140 2917.600 3407.500 ;
        RECT 2.400 3343.540 2917.600 3406.140 ;
        RECT 2.800 3341.540 2917.200 3343.540 ;
        RECT 2.400 3278.940 2917.600 3341.540 ;
        RECT 2.800 3277.580 2917.600 3278.940 ;
        RECT 2.800 3276.940 2917.200 3277.580 ;
        RECT 2.400 3275.580 2917.200 3276.940 ;
        RECT 2.400 3214.340 2917.600 3275.580 ;
        RECT 2.800 3212.340 2917.600 3214.340 ;
        RECT 2.400 3211.620 2917.600 3212.340 ;
        RECT 2.400 3209.620 2917.200 3211.620 ;
        RECT 2.400 3149.740 2917.600 3209.620 ;
        RECT 2.800 3147.740 2917.600 3149.740 ;
        RECT 2.400 3145.660 2917.600 3147.740 ;
        RECT 2.400 3143.660 2917.200 3145.660 ;
        RECT 2.400 3085.140 2917.600 3143.660 ;
        RECT 2.800 3083.140 2917.600 3085.140 ;
        RECT 2.400 3079.700 2917.600 3083.140 ;
        RECT 2.400 3077.700 2917.200 3079.700 ;
        RECT 2.400 3020.540 2917.600 3077.700 ;
        RECT 2.800 3018.540 2917.600 3020.540 ;
        RECT 2.400 3013.740 2917.600 3018.540 ;
        RECT 2.400 3011.740 2917.200 3013.740 ;
        RECT 2.400 2955.940 2917.600 3011.740 ;
        RECT 2.800 2953.940 2917.600 2955.940 ;
        RECT 2.400 2947.780 2917.600 2953.940 ;
        RECT 2.400 2945.780 2917.200 2947.780 ;
        RECT 2.400 2891.340 2917.600 2945.780 ;
        RECT 2.800 2889.340 2917.600 2891.340 ;
        RECT 2.400 2881.820 2917.600 2889.340 ;
        RECT 2.400 2879.820 2917.200 2881.820 ;
        RECT 2.400 2826.740 2917.600 2879.820 ;
        RECT 2.800 2824.740 2917.600 2826.740 ;
        RECT 2.400 2815.860 2917.600 2824.740 ;
        RECT 2.400 2813.860 2917.200 2815.860 ;
        RECT 2.400 2762.140 2917.600 2813.860 ;
        RECT 2.800 2760.140 2917.600 2762.140 ;
        RECT 2.400 2749.900 2917.600 2760.140 ;
        RECT 2.400 2747.900 2917.200 2749.900 ;
        RECT 2.400 2697.540 2917.600 2747.900 ;
        RECT 2.800 2695.540 2917.600 2697.540 ;
        RECT 2.400 2683.940 2917.600 2695.540 ;
        RECT 2.400 2681.940 2917.200 2683.940 ;
        RECT 2.400 2632.940 2917.600 2681.940 ;
        RECT 2.800 2630.940 2917.600 2632.940 ;
        RECT 2.400 2617.980 2917.600 2630.940 ;
        RECT 2.400 2615.980 2917.200 2617.980 ;
        RECT 2.400 2568.340 2917.600 2615.980 ;
        RECT 2.800 2566.340 2917.600 2568.340 ;
        RECT 2.400 2552.020 2917.600 2566.340 ;
        RECT 2.400 2550.020 2917.200 2552.020 ;
        RECT 2.400 2503.740 2917.600 2550.020 ;
        RECT 2.800 2501.740 2917.600 2503.740 ;
        RECT 2.400 2486.060 2917.600 2501.740 ;
        RECT 2.400 2484.060 2917.200 2486.060 ;
        RECT 2.400 2439.140 2917.600 2484.060 ;
        RECT 2.800 2437.140 2917.600 2439.140 ;
        RECT 2.400 2420.100 2917.600 2437.140 ;
        RECT 2.400 2418.100 2917.200 2420.100 ;
        RECT 2.400 2374.540 2917.600 2418.100 ;
        RECT 2.800 2372.540 2917.600 2374.540 ;
        RECT 2.400 2354.140 2917.600 2372.540 ;
        RECT 2.400 2352.140 2917.200 2354.140 ;
        RECT 2.400 2309.940 2917.600 2352.140 ;
        RECT 2.800 2307.940 2917.600 2309.940 ;
        RECT 2.400 2288.180 2917.600 2307.940 ;
        RECT 2.400 2286.180 2917.200 2288.180 ;
        RECT 2.400 2245.340 2917.600 2286.180 ;
        RECT 2.800 2243.340 2917.600 2245.340 ;
        RECT 2.400 2222.220 2917.600 2243.340 ;
        RECT 2.400 2220.220 2917.200 2222.220 ;
        RECT 2.400 2180.740 2917.600 2220.220 ;
        RECT 2.800 2178.740 2917.600 2180.740 ;
        RECT 2.400 2156.260 2917.600 2178.740 ;
        RECT 2.400 2154.260 2917.200 2156.260 ;
        RECT 2.400 2116.140 2917.600 2154.260 ;
        RECT 2.800 2114.140 2917.600 2116.140 ;
        RECT 2.400 2090.300 2917.600 2114.140 ;
        RECT 2.400 2088.300 2917.200 2090.300 ;
        RECT 2.400 2051.540 2917.600 2088.300 ;
        RECT 2.800 2049.540 2917.600 2051.540 ;
        RECT 2.400 2024.340 2917.600 2049.540 ;
        RECT 2.400 2022.340 2917.200 2024.340 ;
        RECT 2.400 1986.940 2917.600 2022.340 ;
        RECT 2.800 1984.940 2917.600 1986.940 ;
        RECT 2.400 1958.380 2917.600 1984.940 ;
        RECT 2.400 1956.380 2917.200 1958.380 ;
        RECT 2.400 1922.340 2917.600 1956.380 ;
        RECT 2.800 1920.340 2917.600 1922.340 ;
        RECT 2.400 1892.420 2917.600 1920.340 ;
        RECT 2.400 1890.420 2917.200 1892.420 ;
        RECT 2.400 1857.740 2917.600 1890.420 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1728.540 2917.600 1758.500 ;
        RECT 2.800 1726.540 2917.600 1728.540 ;
        RECT 2.400 1694.540 2917.600 1726.540 ;
        RECT 2.400 1692.540 2917.200 1694.540 ;
        RECT 2.400 1663.940 2917.600 1692.540 ;
        RECT 2.800 1661.940 2917.600 1663.940 ;
        RECT 2.400 1628.580 2917.600 1661.940 ;
        RECT 2.400 1626.580 2917.200 1628.580 ;
        RECT 2.400 1599.340 2917.600 1626.580 ;
        RECT 2.800 1597.340 2917.600 1599.340 ;
        RECT 2.400 1562.620 2917.600 1597.340 ;
        RECT 2.400 1560.620 2917.200 1562.620 ;
        RECT 2.400 1534.740 2917.600 1560.620 ;
        RECT 2.800 1532.740 2917.600 1534.740 ;
        RECT 2.400 1496.660 2917.600 1532.740 ;
        RECT 2.400 1494.660 2917.200 1496.660 ;
        RECT 2.400 1470.140 2917.600 1494.660 ;
        RECT 2.800 1468.140 2917.600 1470.140 ;
        RECT 2.400 1430.700 2917.600 1468.140 ;
        RECT 2.400 1428.700 2917.200 1430.700 ;
        RECT 2.400 1405.540 2917.600 1428.700 ;
        RECT 2.800 1403.540 2917.600 1405.540 ;
        RECT 2.400 1364.740 2917.600 1403.540 ;
        RECT 2.400 1362.740 2917.200 1364.740 ;
        RECT 2.400 1340.940 2917.600 1362.740 ;
        RECT 2.800 1338.940 2917.600 1340.940 ;
        RECT 2.400 1298.780 2917.600 1338.940 ;
        RECT 2.400 1296.780 2917.200 1298.780 ;
        RECT 2.400 1276.340 2917.600 1296.780 ;
        RECT 2.800 1274.340 2917.600 1276.340 ;
        RECT 2.400 1232.820 2917.600 1274.340 ;
        RECT 2.400 1230.820 2917.200 1232.820 ;
        RECT 2.400 1211.740 2917.600 1230.820 ;
        RECT 2.800 1209.740 2917.600 1211.740 ;
        RECT 2.400 1166.860 2917.600 1209.740 ;
        RECT 2.400 1164.860 2917.200 1166.860 ;
        RECT 2.400 1147.140 2917.600 1164.860 ;
        RECT 2.800 1145.140 2917.600 1147.140 ;
        RECT 2.400 1100.900 2917.600 1145.140 ;
        RECT 2.400 1098.900 2917.200 1100.900 ;
        RECT 2.400 1082.540 2917.600 1098.900 ;
        RECT 2.800 1080.540 2917.600 1082.540 ;
        RECT 2.400 1034.940 2917.600 1080.540 ;
        RECT 2.400 1032.940 2917.200 1034.940 ;
        RECT 2.400 1017.940 2917.600 1032.940 ;
        RECT 2.800 1015.940 2917.600 1017.940 ;
        RECT 2.400 968.980 2917.600 1015.940 ;
        RECT 2.400 966.980 2917.200 968.980 ;
        RECT 2.400 953.340 2917.600 966.980 ;
        RECT 2.800 951.340 2917.600 953.340 ;
        RECT 2.400 903.020 2917.600 951.340 ;
        RECT 2.400 901.020 2917.200 903.020 ;
        RECT 2.400 888.740 2917.600 901.020 ;
        RECT 2.800 886.740 2917.600 888.740 ;
        RECT 2.400 837.060 2917.600 886.740 ;
        RECT 2.400 835.060 2917.200 837.060 ;
        RECT 2.400 824.140 2917.600 835.060 ;
        RECT 2.800 822.140 2917.600 824.140 ;
        RECT 2.400 771.100 2917.600 822.140 ;
        RECT 2.400 769.100 2917.200 771.100 ;
        RECT 2.400 759.540 2917.600 769.100 ;
        RECT 2.800 757.540 2917.600 759.540 ;
        RECT 2.400 705.140 2917.600 757.540 ;
        RECT 2.400 703.140 2917.200 705.140 ;
        RECT 2.400 694.940 2917.600 703.140 ;
        RECT 2.800 692.940 2917.600 694.940 ;
        RECT 2.400 639.180 2917.600 692.940 ;
        RECT 2.400 637.180 2917.200 639.180 ;
        RECT 2.400 630.340 2917.600 637.180 ;
        RECT 2.800 628.340 2917.600 630.340 ;
        RECT 2.400 573.220 2917.600 628.340 ;
        RECT 2.400 571.220 2917.200 573.220 ;
        RECT 2.400 565.740 2917.600 571.220 ;
        RECT 2.800 563.740 2917.600 565.740 ;
        RECT 2.400 507.260 2917.600 563.740 ;
        RECT 2.400 505.260 2917.200 507.260 ;
        RECT 2.400 501.140 2917.600 505.260 ;
        RECT 2.800 499.140 2917.600 501.140 ;
        RECT 2.400 441.300 2917.600 499.140 ;
        RECT 2.400 439.300 2917.200 441.300 ;
        RECT 2.400 436.540 2917.600 439.300 ;
        RECT 2.800 434.540 2917.600 436.540 ;
        RECT 2.400 375.340 2917.600 434.540 ;
        RECT 2.400 373.340 2917.200 375.340 ;
        RECT 2.400 371.940 2917.600 373.340 ;
        RECT 2.800 369.940 2917.600 371.940 ;
        RECT 2.400 309.380 2917.600 369.940 ;
        RECT 2.400 307.380 2917.200 309.380 ;
        RECT 2.400 307.340 2917.600 307.380 ;
        RECT 2.800 305.340 2917.600 307.340 ;
        RECT 2.400 243.420 2917.600 305.340 ;
        RECT 2.400 242.740 2917.200 243.420 ;
        RECT 2.800 241.420 2917.200 242.740 ;
        RECT 2.800 240.740 2917.600 241.420 ;
        RECT 2.400 178.140 2917.600 240.740 ;
        RECT 2.800 177.460 2917.600 178.140 ;
        RECT 2.800 176.140 2917.200 177.460 ;
        RECT 2.400 175.460 2917.200 176.140 ;
        RECT 2.400 113.540 2917.600 175.460 ;
        RECT 2.800 111.540 2917.600 113.540 ;
        RECT 2.400 111.500 2917.600 111.540 ;
        RECT 2.400 109.500 2917.200 111.500 ;
        RECT 2.400 48.940 2917.600 109.500 ;
        RECT 2.800 46.940 2917.600 48.940 ;
        RECT 2.400 45.540 2917.600 46.940 ;
        RECT 2.400 43.540 2917.200 45.540 ;
        RECT 2.400 10.715 2917.600 43.540 ;
      LAYER met4 ;
        RECT 38.935 12.415 39.770 3447.425 ;
        RECT 43.670 12.415 47.870 3447.425 ;
        RECT 51.770 3439.900 123.570 3447.425 ;
        RECT 127.470 3439.900 131.670 3447.425 ;
        RECT 135.570 3439.900 139.770 3447.425 ;
        RECT 143.670 3439.900 147.870 3447.425 ;
        RECT 151.770 3439.900 223.570 3447.425 ;
        RECT 227.470 3439.900 231.670 3447.425 ;
        RECT 235.570 3439.900 239.770 3447.425 ;
        RECT 243.670 3439.900 247.870 3447.425 ;
        RECT 251.770 3439.900 323.570 3447.425 ;
        RECT 327.470 3439.900 331.670 3447.425 ;
        RECT 335.570 3439.900 339.770 3447.425 ;
        RECT 343.670 3439.900 347.870 3447.425 ;
        RECT 351.770 3439.900 423.570 3447.425 ;
        RECT 427.470 3439.900 431.670 3447.425 ;
        RECT 435.570 3439.900 439.770 3447.425 ;
        RECT 443.670 3439.900 447.870 3447.425 ;
        RECT 451.770 3439.900 523.570 3447.425 ;
        RECT 527.470 3439.900 531.670 3447.425 ;
        RECT 535.570 3439.900 539.770 3447.425 ;
        RECT 543.670 3439.900 547.870 3447.425 ;
        RECT 551.770 3439.900 623.570 3447.425 ;
        RECT 627.470 3439.900 631.670 3447.425 ;
        RECT 635.570 3439.900 639.770 3447.425 ;
        RECT 643.670 3439.900 647.870 3447.425 ;
        RECT 651.770 3439.900 723.570 3447.425 ;
        RECT 727.470 3439.900 731.670 3447.425 ;
        RECT 735.570 3439.900 739.770 3447.425 ;
        RECT 743.670 3439.900 747.870 3447.425 ;
        RECT 751.770 3439.900 823.570 3447.425 ;
        RECT 827.470 3439.900 831.670 3447.425 ;
        RECT 835.570 3439.900 839.770 3447.425 ;
        RECT 843.670 3439.900 847.870 3447.425 ;
        RECT 851.770 3439.900 923.570 3447.425 ;
        RECT 927.470 3439.900 931.670 3447.425 ;
        RECT 935.570 3439.900 939.770 3447.425 ;
        RECT 943.670 3439.900 947.870 3447.425 ;
        RECT 951.770 3439.900 1023.570 3447.425 ;
        RECT 1027.470 3439.900 1031.670 3447.425 ;
        RECT 1035.570 3439.900 1039.770 3447.425 ;
        RECT 1043.670 3439.900 1047.870 3447.425 ;
        RECT 1051.770 3439.900 1123.570 3447.425 ;
        RECT 1127.470 3439.900 1131.670 3447.425 ;
        RECT 1135.570 3439.900 1139.770 3447.425 ;
        RECT 1143.670 3439.900 1147.870 3447.425 ;
        RECT 1151.770 3439.900 1223.570 3447.425 ;
        RECT 1227.470 3439.900 1231.670 3447.425 ;
        RECT 1235.570 3439.900 1239.770 3447.425 ;
        RECT 1243.670 3439.900 1247.870 3447.425 ;
        RECT 1251.770 3439.900 1323.570 3447.425 ;
        RECT 1327.470 3439.900 1331.670 3447.425 ;
        RECT 1335.570 3439.900 1339.770 3447.425 ;
        RECT 1343.670 3439.900 1347.870 3447.425 ;
        RECT 1351.770 3439.900 1423.570 3447.425 ;
        RECT 51.770 1820.100 1423.570 3439.900 ;
        RECT 51.770 1725.900 123.570 1820.100 ;
        RECT 127.470 1725.900 131.670 1820.100 ;
        RECT 135.570 1725.900 223.570 1820.100 ;
        RECT 227.470 1725.900 231.670 1820.100 ;
        RECT 235.570 1725.900 323.570 1820.100 ;
        RECT 327.470 1725.900 331.670 1820.100 ;
        RECT 335.570 1725.900 423.570 1820.100 ;
        RECT 427.470 1725.900 431.670 1820.100 ;
        RECT 435.570 1725.900 523.570 1820.100 ;
        RECT 527.470 1725.900 531.670 1820.100 ;
        RECT 535.570 1725.900 623.570 1820.100 ;
        RECT 627.470 1725.900 631.670 1820.100 ;
        RECT 635.570 1725.900 723.570 1820.100 ;
        RECT 727.470 1725.900 731.670 1820.100 ;
        RECT 735.570 1725.900 823.570 1820.100 ;
        RECT 827.470 1725.900 831.670 1820.100 ;
        RECT 835.570 1725.900 923.570 1820.100 ;
        RECT 927.470 1725.900 931.670 1820.100 ;
        RECT 935.570 1725.900 1023.570 1820.100 ;
        RECT 1027.470 1725.900 1031.670 1820.100 ;
        RECT 1035.570 1725.900 1123.570 1820.100 ;
        RECT 1127.470 1725.900 1131.670 1820.100 ;
        RECT 1135.570 1725.900 1223.570 1820.100 ;
        RECT 1227.470 1725.900 1231.670 1820.100 ;
        RECT 1235.570 1725.900 1323.570 1820.100 ;
        RECT 1327.470 1725.900 1331.670 1820.100 ;
        RECT 1335.570 1725.900 1423.570 1820.100 ;
        RECT 51.770 106.100 1423.570 1725.900 ;
        RECT 51.770 12.415 123.570 106.100 ;
        RECT 127.470 12.415 131.670 106.100 ;
        RECT 135.570 12.415 139.770 106.100 ;
        RECT 143.670 12.415 147.870 106.100 ;
        RECT 151.770 12.415 223.570 106.100 ;
        RECT 227.470 12.415 231.670 106.100 ;
        RECT 235.570 12.415 239.770 106.100 ;
        RECT 243.670 12.415 247.870 106.100 ;
        RECT 251.770 12.415 323.570 106.100 ;
        RECT 327.470 12.415 331.670 106.100 ;
        RECT 335.570 12.415 339.770 106.100 ;
        RECT 343.670 12.415 347.870 106.100 ;
        RECT 351.770 12.415 423.570 106.100 ;
        RECT 427.470 12.415 431.670 106.100 ;
        RECT 435.570 12.415 439.770 106.100 ;
        RECT 443.670 12.415 447.870 106.100 ;
        RECT 451.770 12.415 523.570 106.100 ;
        RECT 527.470 12.415 531.670 106.100 ;
        RECT 535.570 12.415 539.770 106.100 ;
        RECT 543.670 12.415 547.870 106.100 ;
        RECT 551.770 12.415 623.570 106.100 ;
        RECT 627.470 12.415 631.670 106.100 ;
        RECT 635.570 12.415 639.770 106.100 ;
        RECT 643.670 12.415 647.870 106.100 ;
        RECT 651.770 12.415 723.570 106.100 ;
        RECT 727.470 12.415 731.670 106.100 ;
        RECT 735.570 12.415 739.770 106.100 ;
        RECT 743.670 12.415 747.870 106.100 ;
        RECT 751.770 12.415 823.570 106.100 ;
        RECT 827.470 12.415 831.670 106.100 ;
        RECT 835.570 12.415 839.770 106.100 ;
        RECT 843.670 12.415 847.870 106.100 ;
        RECT 851.770 12.415 923.570 106.100 ;
        RECT 927.470 12.415 931.670 106.100 ;
        RECT 935.570 12.415 939.770 106.100 ;
        RECT 943.670 12.415 947.870 106.100 ;
        RECT 951.770 12.415 1023.570 106.100 ;
        RECT 1027.470 12.415 1031.670 106.100 ;
        RECT 1035.570 12.415 1039.770 106.100 ;
        RECT 1043.670 12.415 1047.870 106.100 ;
        RECT 1051.770 12.415 1123.570 106.100 ;
        RECT 1127.470 12.415 1131.670 106.100 ;
        RECT 1135.570 12.415 1139.770 106.100 ;
        RECT 1143.670 12.415 1147.870 106.100 ;
        RECT 1151.770 12.415 1223.570 106.100 ;
        RECT 1227.470 12.415 1231.670 106.100 ;
        RECT 1235.570 12.415 1239.770 106.100 ;
        RECT 1243.670 12.415 1247.870 106.100 ;
        RECT 1251.770 12.415 1323.570 106.100 ;
        RECT 1327.470 12.415 1331.670 106.100 ;
        RECT 1335.570 12.415 1339.770 106.100 ;
        RECT 1343.670 12.415 1347.870 106.100 ;
        RECT 1351.770 12.415 1423.570 106.100 ;
        RECT 1427.470 12.415 1431.670 3447.425 ;
        RECT 1435.570 12.415 1439.770 3447.425 ;
        RECT 1443.670 12.415 1447.870 3447.425 ;
        RECT 1451.770 3439.900 1523.570 3447.425 ;
        RECT 1527.470 3439.900 1531.670 3447.425 ;
        RECT 1535.570 3439.900 1539.770 3447.425 ;
        RECT 1543.670 3439.900 1547.870 3447.425 ;
        RECT 1551.770 3439.900 1623.570 3447.425 ;
        RECT 1627.470 3439.900 1631.670 3447.425 ;
        RECT 1635.570 3439.900 1639.770 3447.425 ;
        RECT 1643.670 3439.900 1647.870 3447.425 ;
        RECT 1651.770 3439.900 1723.570 3447.425 ;
        RECT 1727.470 3439.900 1731.670 3447.425 ;
        RECT 1735.570 3439.900 1739.770 3447.425 ;
        RECT 1743.670 3439.900 1747.870 3447.425 ;
        RECT 1751.770 3439.900 1823.570 3447.425 ;
        RECT 1827.470 3439.900 1831.670 3447.425 ;
        RECT 1835.570 3439.900 1839.770 3447.425 ;
        RECT 1843.670 3439.900 1847.870 3447.425 ;
        RECT 1851.770 3439.900 1923.570 3447.425 ;
        RECT 1927.470 3439.900 1931.670 3447.425 ;
        RECT 1935.570 3439.900 1939.770 3447.425 ;
        RECT 1943.670 3439.900 1947.870 3447.425 ;
        RECT 1951.770 3439.900 2023.570 3447.425 ;
        RECT 2027.470 3439.900 2031.670 3447.425 ;
        RECT 2035.570 3439.900 2039.770 3447.425 ;
        RECT 2043.670 3439.900 2047.870 3447.425 ;
        RECT 2051.770 3439.900 2123.570 3447.425 ;
        RECT 2127.470 3439.900 2131.670 3447.425 ;
        RECT 2135.570 3439.900 2139.770 3447.425 ;
        RECT 2143.670 3439.900 2147.870 3447.425 ;
        RECT 2151.770 3439.900 2223.570 3447.425 ;
        RECT 2227.470 3439.900 2231.670 3447.425 ;
        RECT 2235.570 3439.900 2239.770 3447.425 ;
        RECT 2243.670 3439.900 2247.870 3447.425 ;
        RECT 2251.770 3439.900 2323.570 3447.425 ;
        RECT 2327.470 3439.900 2331.670 3447.425 ;
        RECT 2335.570 3439.900 2339.770 3447.425 ;
        RECT 2343.670 3439.900 2347.870 3447.425 ;
        RECT 2351.770 3439.900 2423.570 3447.425 ;
        RECT 2427.470 3439.900 2431.670 3447.425 ;
        RECT 2435.570 3439.900 2439.770 3447.425 ;
        RECT 2443.670 3439.900 2447.870 3447.425 ;
        RECT 2451.770 3439.900 2523.570 3447.425 ;
        RECT 2527.470 3439.900 2531.670 3447.425 ;
        RECT 2535.570 3439.900 2539.770 3447.425 ;
        RECT 2543.670 3439.900 2547.870 3447.425 ;
        RECT 2551.770 3439.900 2623.570 3447.425 ;
        RECT 2627.470 3439.900 2631.670 3447.425 ;
        RECT 2635.570 3439.900 2639.770 3447.425 ;
        RECT 2643.670 3439.900 2647.870 3447.425 ;
        RECT 2651.770 3439.900 2723.570 3447.425 ;
        RECT 2727.470 3439.900 2731.670 3447.425 ;
        RECT 2735.570 3439.900 2739.770 3447.425 ;
        RECT 2743.670 3439.900 2747.870 3447.425 ;
        RECT 2751.770 3439.900 2823.570 3447.425 ;
        RECT 2827.470 3439.900 2831.670 3447.425 ;
        RECT 2835.570 3439.900 2839.770 3447.425 ;
        RECT 2843.670 3439.900 2847.870 3447.425 ;
        RECT 1451.770 1820.100 2847.870 3439.900 ;
        RECT 1451.770 1725.900 1523.570 1820.100 ;
        RECT 1527.470 1725.900 1531.670 1820.100 ;
        RECT 1535.570 1725.900 1623.570 1820.100 ;
        RECT 1627.470 1725.900 1631.670 1820.100 ;
        RECT 1635.570 1725.900 1723.570 1820.100 ;
        RECT 1727.470 1725.900 1731.670 1820.100 ;
        RECT 1735.570 1725.900 1823.570 1820.100 ;
        RECT 1827.470 1725.900 1831.670 1820.100 ;
        RECT 1835.570 1725.900 1923.570 1820.100 ;
        RECT 1927.470 1725.900 1931.670 1820.100 ;
        RECT 1935.570 1725.900 2023.570 1820.100 ;
        RECT 2027.470 1725.900 2031.670 1820.100 ;
        RECT 2035.570 1725.900 2123.570 1820.100 ;
        RECT 2127.470 1725.900 2131.670 1820.100 ;
        RECT 2135.570 1725.900 2223.570 1820.100 ;
        RECT 2227.470 1725.900 2231.670 1820.100 ;
        RECT 2235.570 1725.900 2323.570 1820.100 ;
        RECT 2327.470 1725.900 2331.670 1820.100 ;
        RECT 2335.570 1725.900 2423.570 1820.100 ;
        RECT 2427.470 1725.900 2431.670 1820.100 ;
        RECT 2435.570 1725.900 2523.570 1820.100 ;
        RECT 2527.470 1725.900 2531.670 1820.100 ;
        RECT 2535.570 1725.900 2623.570 1820.100 ;
        RECT 2627.470 1725.900 2631.670 1820.100 ;
        RECT 2635.570 1725.900 2723.570 1820.100 ;
        RECT 2727.470 1725.900 2731.670 1820.100 ;
        RECT 2735.570 1725.900 2823.570 1820.100 ;
        RECT 2827.470 1725.900 2831.670 1820.100 ;
        RECT 2835.570 1725.900 2847.870 1820.100 ;
        RECT 1451.770 106.100 2847.870 1725.900 ;
        RECT 1451.770 12.415 1523.570 106.100 ;
        RECT 1527.470 12.415 1531.670 106.100 ;
        RECT 1535.570 12.415 1539.770 106.100 ;
        RECT 1543.670 12.415 1547.870 106.100 ;
        RECT 1551.770 12.415 1623.570 106.100 ;
        RECT 1627.470 12.415 1631.670 106.100 ;
        RECT 1635.570 12.415 1639.770 106.100 ;
        RECT 1643.670 12.415 1647.870 106.100 ;
        RECT 1651.770 12.415 1723.570 106.100 ;
        RECT 1727.470 12.415 1731.670 106.100 ;
        RECT 1735.570 12.415 1739.770 106.100 ;
        RECT 1743.670 12.415 1747.870 106.100 ;
        RECT 1751.770 12.415 1823.570 106.100 ;
        RECT 1827.470 12.415 1831.670 106.100 ;
        RECT 1835.570 12.415 1839.770 106.100 ;
        RECT 1843.670 12.415 1847.870 106.100 ;
        RECT 1851.770 12.415 1923.570 106.100 ;
        RECT 1927.470 12.415 1931.670 106.100 ;
        RECT 1935.570 12.415 1939.770 106.100 ;
        RECT 1943.670 12.415 1947.870 106.100 ;
        RECT 1951.770 12.415 2023.570 106.100 ;
        RECT 2027.470 12.415 2031.670 106.100 ;
        RECT 2035.570 12.415 2039.770 106.100 ;
        RECT 2043.670 12.415 2047.870 106.100 ;
        RECT 2051.770 12.415 2123.570 106.100 ;
        RECT 2127.470 12.415 2131.670 106.100 ;
        RECT 2135.570 12.415 2139.770 106.100 ;
        RECT 2143.670 12.415 2147.870 106.100 ;
        RECT 2151.770 12.415 2223.570 106.100 ;
        RECT 2227.470 12.415 2231.670 106.100 ;
        RECT 2235.570 12.415 2239.770 106.100 ;
        RECT 2243.670 12.415 2247.870 106.100 ;
        RECT 2251.770 12.415 2323.570 106.100 ;
        RECT 2327.470 12.415 2331.670 106.100 ;
        RECT 2335.570 12.415 2339.770 106.100 ;
        RECT 2343.670 12.415 2347.870 106.100 ;
        RECT 2351.770 12.415 2423.570 106.100 ;
        RECT 2427.470 12.415 2431.670 106.100 ;
        RECT 2435.570 12.415 2439.770 106.100 ;
        RECT 2443.670 12.415 2447.870 106.100 ;
        RECT 2451.770 12.415 2523.570 106.100 ;
        RECT 2527.470 12.415 2531.670 106.100 ;
        RECT 2535.570 12.415 2539.770 106.100 ;
        RECT 2543.670 12.415 2547.870 106.100 ;
        RECT 2551.770 12.415 2623.570 106.100 ;
        RECT 2627.470 12.415 2631.670 106.100 ;
        RECT 2635.570 12.415 2639.770 106.100 ;
        RECT 2643.670 12.415 2647.870 106.100 ;
        RECT 2651.770 12.415 2723.570 106.100 ;
        RECT 2727.470 12.415 2731.670 106.100 ;
        RECT 2735.570 12.415 2739.770 106.100 ;
        RECT 2743.670 12.415 2747.870 106.100 ;
        RECT 2751.770 12.415 2823.570 106.100 ;
        RECT 2827.470 12.415 2831.670 106.100 ;
        RECT 2835.570 12.415 2839.770 106.100 ;
        RECT 2843.670 12.415 2847.870 106.100 ;
        RECT 2851.770 12.415 2871.945 3447.425 ;
      LAYER met5 ;
        RECT 559.940 1658.330 1784.220 1726.300 ;
        RECT 559.940 1650.230 1784.220 1652.030 ;
        RECT 559.940 1642.130 1784.220 1643.930 ;
        RECT 559.940 1634.030 1784.220 1635.830 ;
        RECT 559.940 1558.330 1784.220 1627.730 ;
        RECT 559.940 1550.230 1784.220 1552.030 ;
        RECT 559.940 1542.130 1784.220 1543.930 ;
        RECT 559.940 1534.030 1784.220 1535.830 ;
        RECT 559.940 1458.330 1784.220 1527.730 ;
        RECT 559.940 1450.230 1784.220 1452.030 ;
        RECT 559.940 1442.130 1784.220 1443.930 ;
        RECT 559.940 1434.030 1784.220 1435.830 ;
        RECT 559.940 1358.330 1784.220 1427.730 ;
        RECT 559.940 1350.230 1784.220 1352.030 ;
        RECT 559.940 1342.130 1784.220 1343.930 ;
        RECT 559.940 1334.030 1784.220 1335.830 ;
        RECT 559.940 1258.330 1784.220 1327.730 ;
        RECT 559.940 1250.230 1784.220 1252.030 ;
        RECT 559.940 1242.130 1784.220 1243.930 ;
        RECT 559.940 1234.030 1784.220 1235.830 ;
        RECT 559.940 1158.330 1784.220 1227.730 ;
        RECT 559.940 1150.230 1784.220 1152.030 ;
        RECT 559.940 1142.130 1784.220 1143.930 ;
        RECT 559.940 1134.030 1784.220 1135.830 ;
        RECT 559.940 1058.330 1784.220 1127.730 ;
        RECT 559.940 1050.230 1784.220 1052.030 ;
        RECT 559.940 1042.130 1784.220 1043.930 ;
        RECT 559.940 1034.030 1784.220 1035.830 ;
        RECT 559.940 958.330 1784.220 1027.730 ;
        RECT 559.940 950.230 1784.220 952.030 ;
        RECT 559.940 942.130 1784.220 943.930 ;
        RECT 559.940 934.030 1784.220 935.830 ;
        RECT 559.940 858.330 1784.220 927.730 ;
        RECT 559.940 850.230 1784.220 852.030 ;
        RECT 559.940 842.130 1784.220 843.930 ;
        RECT 559.940 834.030 1784.220 835.830 ;
        RECT 559.940 758.330 1784.220 827.730 ;
        RECT 559.940 750.230 1784.220 752.030 ;
        RECT 559.940 742.130 1784.220 743.930 ;
        RECT 559.940 734.030 1784.220 735.830 ;
        RECT 559.940 658.330 1784.220 727.730 ;
        RECT 559.940 650.230 1784.220 652.030 ;
        RECT 559.940 642.130 1784.220 643.930 ;
        RECT 559.940 634.030 1784.220 635.830 ;
        RECT 559.940 558.330 1784.220 627.730 ;
        RECT 559.940 550.230 1784.220 552.030 ;
        RECT 559.940 542.130 1784.220 543.930 ;
        RECT 559.940 534.030 1784.220 535.830 ;
        RECT 559.940 458.330 1784.220 527.730 ;
        RECT 559.940 450.230 1784.220 452.030 ;
        RECT 559.940 442.130 1784.220 443.930 ;
        RECT 559.940 434.030 1784.220 435.830 ;
        RECT 559.940 358.330 1784.220 427.730 ;
        RECT 559.940 350.230 1784.220 352.030 ;
        RECT 559.940 342.130 1784.220 343.930 ;
        RECT 559.940 334.030 1784.220 335.830 ;
        RECT 559.940 258.330 1784.220 327.730 ;
        RECT 559.940 250.230 1784.220 252.030 ;
        RECT 559.940 242.130 1784.220 243.930 ;
        RECT 559.940 234.030 1784.220 235.830 ;
        RECT 559.940 158.330 1784.220 227.730 ;
        RECT 559.940 150.230 1784.220 152.030 ;
        RECT 559.940 142.130 1784.220 143.930 ;
        RECT 559.940 134.030 1784.220 135.830 ;
        RECT 559.940 58.700 1784.220 127.730 ;
  END
END user_project_wrapper
END LIBRARY

