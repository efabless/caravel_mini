magic
tech sky130A
magscale 1 2
timestamp 1682300533
<< obsli1 >>
rect 1104 2159 258888 317713
<< obsm1 >>
rect 1104 1640 259058 317892
<< metal2 >>
rect 5510 319520 5622 320960
rect 15078 319520 15190 320960
rect 24646 319520 24758 320960
rect 34214 319520 34326 320960
rect 43782 319520 43894 320960
rect 53350 319520 53462 320960
rect 62918 319520 63030 320960
rect 72486 319520 72598 320960
rect 82054 319520 82166 320960
rect 91622 319520 91734 320960
rect 101190 319520 101302 320960
rect 110758 319520 110870 320960
rect 120326 319520 120438 320960
rect 129894 319520 130006 320960
rect 139462 319520 139574 320960
rect 149030 319520 149142 320960
rect 158598 319520 158710 320960
rect 168166 319520 168278 320960
rect 177734 319520 177846 320960
rect 187302 319520 187414 320960
rect 196870 319520 196982 320960
rect 206438 319520 206550 320960
rect 216006 319520 216118 320960
rect 225574 319520 225686 320960
rect 235142 319520 235254 320960
rect 244710 319520 244822 320960
rect 254278 319520 254390 320960
rect 6706 -960 6818 480
rect 8454 -960 8566 480
rect 10202 -960 10314 480
rect 11950 -960 12062 480
rect 13698 -960 13810 480
rect 15446 -960 15558 480
rect 17194 -960 17306 480
rect 18942 -960 19054 480
rect 20690 -960 20802 480
rect 22438 -960 22550 480
rect 24186 -960 24298 480
rect 25934 -960 26046 480
rect 27682 -960 27794 480
rect 29430 -960 29542 480
rect 31178 -960 31290 480
rect 32926 -960 33038 480
rect 34674 -960 34786 480
rect 36422 -960 36534 480
rect 38170 -960 38282 480
rect 39918 -960 40030 480
rect 41666 -960 41778 480
rect 43414 -960 43526 480
rect 45162 -960 45274 480
rect 46910 -960 47022 480
rect 48658 -960 48770 480
rect 50406 -960 50518 480
rect 52154 -960 52266 480
rect 53902 -960 54014 480
rect 55650 -960 55762 480
rect 57398 -960 57510 480
rect 59146 -960 59258 480
rect 60894 -960 61006 480
rect 62642 -960 62754 480
rect 64390 -960 64502 480
rect 66138 -960 66250 480
rect 67886 -960 67998 480
rect 69634 -960 69746 480
rect 71382 -960 71494 480
rect 73130 -960 73242 480
rect 74878 -960 74990 480
rect 76626 -960 76738 480
rect 78374 -960 78486 480
rect 80122 -960 80234 480
rect 81870 -960 81982 480
rect 83618 -960 83730 480
rect 85366 -960 85478 480
rect 87114 -960 87226 480
rect 88862 -960 88974 480
rect 90610 -960 90722 480
rect 92358 -960 92470 480
rect 94106 -960 94218 480
rect 95854 -960 95966 480
rect 97602 -960 97714 480
rect 99350 -960 99462 480
rect 101098 -960 101210 480
rect 102846 -960 102958 480
rect 104594 -960 104706 480
rect 106342 -960 106454 480
rect 108090 -960 108202 480
rect 109838 -960 109950 480
rect 111586 -960 111698 480
rect 113334 -960 113446 480
rect 115082 -960 115194 480
rect 116830 -960 116942 480
rect 118578 -960 118690 480
rect 120326 -960 120438 480
rect 122074 -960 122186 480
rect 123822 -960 123934 480
rect 125570 -960 125682 480
rect 127318 -960 127430 480
rect 129066 -960 129178 480
rect 130814 -960 130926 480
rect 132562 -960 132674 480
rect 134310 -960 134422 480
rect 136058 -960 136170 480
rect 137806 -960 137918 480
rect 139554 -960 139666 480
rect 141302 -960 141414 480
rect 143050 -960 143162 480
rect 144798 -960 144910 480
rect 146546 -960 146658 480
rect 148294 -960 148406 480
rect 150042 -960 150154 480
rect 151790 -960 151902 480
rect 153538 -960 153650 480
rect 155286 -960 155398 480
rect 157034 -960 157146 480
rect 158782 -960 158894 480
rect 160530 -960 160642 480
rect 162278 -960 162390 480
rect 164026 -960 164138 480
rect 165774 -960 165886 480
rect 167522 -960 167634 480
rect 169270 -960 169382 480
rect 171018 -960 171130 480
rect 172766 -960 172878 480
rect 174514 -960 174626 480
rect 176262 -960 176374 480
rect 178010 -960 178122 480
rect 179758 -960 179870 480
rect 181506 -960 181618 480
rect 183254 -960 183366 480
rect 185002 -960 185114 480
rect 186750 -960 186862 480
rect 188498 -960 188610 480
rect 190246 -960 190358 480
rect 191994 -960 192106 480
rect 193742 -960 193854 480
rect 195490 -960 195602 480
rect 197238 -960 197350 480
rect 198986 -960 199098 480
rect 200734 -960 200846 480
rect 202482 -960 202594 480
rect 204230 -960 204342 480
rect 205978 -960 206090 480
rect 207726 -960 207838 480
rect 209474 -960 209586 480
rect 211222 -960 211334 480
rect 212970 -960 213082 480
rect 214718 -960 214830 480
rect 216466 -960 216578 480
rect 218214 -960 218326 480
rect 219962 -960 220074 480
rect 221710 -960 221822 480
rect 223458 -960 223570 480
rect 225206 -960 225318 480
rect 226954 -960 227066 480
rect 228702 -960 228814 480
rect 230450 -960 230562 480
rect 232198 -960 232310 480
rect 233946 -960 234058 480
rect 235694 -960 235806 480
rect 237442 -960 237554 480
rect 239190 -960 239302 480
rect 240938 -960 241050 480
rect 242686 -960 242798 480
rect 244434 -960 244546 480
rect 246182 -960 246294 480
rect 247930 -960 248042 480
rect 249678 -960 249790 480
rect 251426 -960 251538 480
rect 253174 -960 253286 480
<< obsm2 >>
rect 1398 319464 5454 319520
rect 5678 319464 15022 319520
rect 15246 319464 24590 319520
rect 24814 319464 34158 319520
rect 34382 319464 43726 319520
rect 43950 319464 53294 319520
rect 53518 319464 62862 319520
rect 63086 319464 72430 319520
rect 72654 319464 81998 319520
rect 82222 319464 91566 319520
rect 91790 319464 101134 319520
rect 101358 319464 110702 319520
rect 110926 319464 120270 319520
rect 120494 319464 129838 319520
rect 130062 319464 139406 319520
rect 139630 319464 148974 319520
rect 149198 319464 158542 319520
rect 158766 319464 168110 319520
rect 168334 319464 177678 319520
rect 177902 319464 187246 319520
rect 187470 319464 196814 319520
rect 197038 319464 206382 319520
rect 206606 319464 215950 319520
rect 216174 319464 225518 319520
rect 225742 319464 235086 319520
rect 235310 319464 244654 319520
rect 244878 319464 254222 319520
rect 254446 319464 259052 319520
rect 1398 536 259052 319464
rect 1398 326 6650 536
rect 6874 326 8398 536
rect 8622 326 10146 536
rect 10370 326 11894 536
rect 12118 326 13642 536
rect 13866 326 15390 536
rect 15614 326 17138 536
rect 17362 326 18886 536
rect 19110 326 20634 536
rect 20858 326 22382 536
rect 22606 326 24130 536
rect 24354 326 25878 536
rect 26102 326 27626 536
rect 27850 326 29374 536
rect 29598 326 31122 536
rect 31346 326 32870 536
rect 33094 326 34618 536
rect 34842 326 36366 536
rect 36590 326 38114 536
rect 38338 326 39862 536
rect 40086 326 41610 536
rect 41834 326 43358 536
rect 43582 326 45106 536
rect 45330 326 46854 536
rect 47078 326 48602 536
rect 48826 326 50350 536
rect 50574 326 52098 536
rect 52322 326 53846 536
rect 54070 326 55594 536
rect 55818 326 57342 536
rect 57566 326 59090 536
rect 59314 326 60838 536
rect 61062 326 62586 536
rect 62810 326 64334 536
rect 64558 326 66082 536
rect 66306 326 67830 536
rect 68054 326 69578 536
rect 69802 326 71326 536
rect 71550 326 73074 536
rect 73298 326 74822 536
rect 75046 326 76570 536
rect 76794 326 78318 536
rect 78542 326 80066 536
rect 80290 326 81814 536
rect 82038 326 83562 536
rect 83786 326 85310 536
rect 85534 326 87058 536
rect 87282 326 88806 536
rect 89030 326 90554 536
rect 90778 326 92302 536
rect 92526 326 94050 536
rect 94274 326 95798 536
rect 96022 326 97546 536
rect 97770 326 99294 536
rect 99518 326 101042 536
rect 101266 326 102790 536
rect 103014 326 104538 536
rect 104762 326 106286 536
rect 106510 326 108034 536
rect 108258 326 109782 536
rect 110006 326 111530 536
rect 111754 326 113278 536
rect 113502 326 115026 536
rect 115250 326 116774 536
rect 116998 326 118522 536
rect 118746 326 120270 536
rect 120494 326 122018 536
rect 122242 326 123766 536
rect 123990 326 125514 536
rect 125738 326 127262 536
rect 127486 326 129010 536
rect 129234 326 130758 536
rect 130982 326 132506 536
rect 132730 326 134254 536
rect 134478 326 136002 536
rect 136226 326 137750 536
rect 137974 326 139498 536
rect 139722 326 141246 536
rect 141470 326 142994 536
rect 143218 326 144742 536
rect 144966 326 146490 536
rect 146714 326 148238 536
rect 148462 326 149986 536
rect 150210 326 151734 536
rect 151958 326 153482 536
rect 153706 326 155230 536
rect 155454 326 156978 536
rect 157202 326 158726 536
rect 158950 326 160474 536
rect 160698 326 162222 536
rect 162446 326 163970 536
rect 164194 326 165718 536
rect 165942 326 167466 536
rect 167690 326 169214 536
rect 169438 326 170962 536
rect 171186 326 172710 536
rect 172934 326 174458 536
rect 174682 326 176206 536
rect 176430 326 177954 536
rect 178178 326 179702 536
rect 179926 326 181450 536
rect 181674 326 183198 536
rect 183422 326 184946 536
rect 185170 326 186694 536
rect 186918 326 188442 536
rect 188666 326 190190 536
rect 190414 326 191938 536
rect 192162 326 193686 536
rect 193910 326 195434 536
rect 195658 326 197182 536
rect 197406 326 198930 536
rect 199154 326 200678 536
rect 200902 326 202426 536
rect 202650 326 204174 536
rect 204398 326 205922 536
rect 206146 326 207670 536
rect 207894 326 209418 536
rect 209642 326 211166 536
rect 211390 326 212914 536
rect 213138 326 214662 536
rect 214886 326 216410 536
rect 216634 326 218158 536
rect 218382 326 219906 536
rect 220130 326 221654 536
rect 221878 326 223402 536
rect 223626 326 225150 536
rect 225374 326 226898 536
rect 227122 326 228646 536
rect 228870 326 230394 536
rect 230618 326 232142 536
rect 232366 326 233890 536
rect 234114 326 235638 536
rect 235862 326 237386 536
rect 237610 326 239134 536
rect 239358 326 240882 536
rect 241106 326 242630 536
rect 242854 326 244378 536
rect 244602 326 246126 536
rect 246350 326 247874 536
rect 248098 326 249622 536
rect 249846 326 251370 536
rect 251594 326 253118 536
rect 253342 326 259052 536
<< metal3 >>
rect -960 314788 480 315028
rect 259520 314924 260960 315164
rect 259520 310844 260960 311084
rect -960 310164 480 310404
rect 259520 306764 260960 307004
rect -960 305540 480 305780
rect 259520 302684 260960 302924
rect -960 300916 480 301156
rect 259520 298604 260960 298844
rect -960 296292 480 296532
rect 259520 294524 260960 294764
rect -960 291668 480 291908
rect 259520 290444 260960 290684
rect -960 287044 480 287284
rect 259520 286364 260960 286604
rect -960 282420 480 282660
rect 259520 282284 260960 282524
rect 259520 278204 260960 278444
rect -960 277796 480 278036
rect 259520 274124 260960 274364
rect -960 273172 480 273412
rect 259520 270044 260960 270284
rect -960 268548 480 268788
rect 259520 265964 260960 266204
rect -960 263924 480 264164
rect 259520 261884 260960 262124
rect -960 259300 480 259540
rect 259520 257804 260960 258044
rect -960 254676 480 254916
rect 259520 253724 260960 253964
rect -960 250052 480 250292
rect 259520 249644 260960 249884
rect -960 245428 480 245668
rect 259520 245564 260960 245804
rect 259520 241484 260960 241724
rect -960 240804 480 241044
rect 259520 237404 260960 237644
rect -960 236180 480 236420
rect 259520 233324 260960 233564
rect -960 231556 480 231796
rect 259520 229244 260960 229484
rect -960 226932 480 227172
rect 259520 225164 260960 225404
rect -960 222308 480 222548
rect 259520 221084 260960 221324
rect -960 217684 480 217924
rect 259520 217004 260960 217244
rect -960 213060 480 213300
rect 259520 212924 260960 213164
rect 259520 208844 260960 209084
rect -960 208436 480 208676
rect 259520 204764 260960 205004
rect -960 203812 480 204052
rect 259520 200684 260960 200924
rect -960 199188 480 199428
rect 259520 196604 260960 196844
rect -960 194564 480 194804
rect 259520 192524 260960 192764
rect -960 189940 480 190180
rect 259520 188444 260960 188684
rect -960 185316 480 185556
rect 259520 184364 260960 184604
rect -960 180692 480 180932
rect 259520 180284 260960 180524
rect -960 176068 480 176308
rect 259520 176204 260960 176444
rect 259520 172124 260960 172364
rect -960 171444 480 171684
rect 259520 168044 260960 168284
rect -960 166820 480 167060
rect 259520 163964 260960 164204
rect -960 162196 480 162436
rect 259520 159884 260960 160124
rect -960 157572 480 157812
rect 259520 155804 260960 156044
rect -960 152948 480 153188
rect 259520 151724 260960 151964
rect -960 148324 480 148564
rect 259520 147644 260960 147884
rect -960 143700 480 143940
rect 259520 143564 260960 143804
rect 259520 139484 260960 139724
rect -960 139076 480 139316
rect 259520 135404 260960 135644
rect -960 134452 480 134692
rect 259520 131324 260960 131564
rect -960 129828 480 130068
rect 259520 127244 260960 127484
rect -960 125204 480 125444
rect 259520 123164 260960 123404
rect -960 120580 480 120820
rect 259520 119084 260960 119324
rect -960 115956 480 116196
rect 259520 115004 260960 115244
rect -960 111332 480 111572
rect 259520 110924 260960 111164
rect -960 106708 480 106948
rect 259520 106844 260960 107084
rect 259520 102764 260960 103004
rect -960 102084 480 102324
rect 259520 98684 260960 98924
rect -960 97460 480 97700
rect 259520 94604 260960 94844
rect -960 92836 480 93076
rect 259520 90524 260960 90764
rect -960 88212 480 88452
rect 259520 86444 260960 86684
rect -960 83588 480 83828
rect 259520 82364 260960 82604
rect -960 78964 480 79204
rect 259520 78284 260960 78524
rect -960 74340 480 74580
rect 259520 74204 260960 74444
rect 259520 70124 260960 70364
rect -960 69716 480 69956
rect 259520 66044 260960 66284
rect -960 65092 480 65332
rect 259520 61964 260960 62204
rect -960 60468 480 60708
rect 259520 57884 260960 58124
rect -960 55844 480 56084
rect 259520 53804 260960 54044
rect -960 51220 480 51460
rect 259520 49724 260960 49964
rect -960 46596 480 46836
rect 259520 45644 260960 45884
rect -960 41972 480 42212
rect 259520 41564 260960 41804
rect -960 37348 480 37588
rect 259520 37484 260960 37724
rect 259520 33404 260960 33644
rect -960 32724 480 32964
rect 259520 29324 260960 29564
rect -960 28100 480 28340
rect 259520 25244 260960 25484
rect -960 23476 480 23716
rect 259520 21164 260960 21404
rect -960 18852 480 19092
rect 259520 17084 260960 17324
rect -960 14228 480 14468
rect 259520 13004 260960 13244
rect -960 9604 480 9844
rect 259520 8924 260960 9164
rect -960 4980 480 5220
rect 259520 4844 260960 5084
<< obsm3 >>
rect 480 315244 259520 317729
rect 480 315108 259440 315244
rect 560 314844 259440 315108
rect 560 314708 259520 314844
rect 480 311164 259520 314708
rect 480 310764 259440 311164
rect 480 310484 259520 310764
rect 560 310084 259520 310484
rect 480 307084 259520 310084
rect 480 306684 259440 307084
rect 480 305860 259520 306684
rect 560 305460 259520 305860
rect 480 303004 259520 305460
rect 480 302604 259440 303004
rect 480 301236 259520 302604
rect 560 300836 259520 301236
rect 480 298924 259520 300836
rect 480 298524 259440 298924
rect 480 296612 259520 298524
rect 560 296212 259520 296612
rect 480 294844 259520 296212
rect 480 294444 259440 294844
rect 480 291988 259520 294444
rect 560 291588 259520 291988
rect 480 290764 259520 291588
rect 480 290364 259440 290764
rect 480 287364 259520 290364
rect 560 286964 259520 287364
rect 480 286684 259520 286964
rect 480 286284 259440 286684
rect 480 282740 259520 286284
rect 560 282604 259520 282740
rect 560 282340 259440 282604
rect 480 282204 259440 282340
rect 480 278524 259520 282204
rect 480 278124 259440 278524
rect 480 278116 259520 278124
rect 560 277716 259520 278116
rect 480 274444 259520 277716
rect 480 274044 259440 274444
rect 480 273492 259520 274044
rect 560 273092 259520 273492
rect 480 270364 259520 273092
rect 480 269964 259440 270364
rect 480 268868 259520 269964
rect 560 268468 259520 268868
rect 480 266284 259520 268468
rect 480 265884 259440 266284
rect 480 264244 259520 265884
rect 560 263844 259520 264244
rect 480 262204 259520 263844
rect 480 261804 259440 262204
rect 480 259620 259520 261804
rect 560 259220 259520 259620
rect 480 258124 259520 259220
rect 480 257724 259440 258124
rect 480 254996 259520 257724
rect 560 254596 259520 254996
rect 480 254044 259520 254596
rect 480 253644 259440 254044
rect 480 250372 259520 253644
rect 560 249972 259520 250372
rect 480 249964 259520 249972
rect 480 249564 259440 249964
rect 480 245884 259520 249564
rect 480 245748 259440 245884
rect 560 245484 259440 245748
rect 560 245348 259520 245484
rect 480 241804 259520 245348
rect 480 241404 259440 241804
rect 480 241124 259520 241404
rect 560 240724 259520 241124
rect 480 237724 259520 240724
rect 480 237324 259440 237724
rect 480 236500 259520 237324
rect 560 236100 259520 236500
rect 480 233644 259520 236100
rect 480 233244 259440 233644
rect 480 231876 259520 233244
rect 560 231476 259520 231876
rect 480 229564 259520 231476
rect 480 229164 259440 229564
rect 480 227252 259520 229164
rect 560 226852 259520 227252
rect 480 225484 259520 226852
rect 480 225084 259440 225484
rect 480 222628 259520 225084
rect 560 222228 259520 222628
rect 480 221404 259520 222228
rect 480 221004 259440 221404
rect 480 218004 259520 221004
rect 560 217604 259520 218004
rect 480 217324 259520 217604
rect 480 216924 259440 217324
rect 480 213380 259520 216924
rect 560 213244 259520 213380
rect 560 212980 259440 213244
rect 480 212844 259440 212980
rect 480 209164 259520 212844
rect 480 208764 259440 209164
rect 480 208756 259520 208764
rect 560 208356 259520 208756
rect 480 205084 259520 208356
rect 480 204684 259440 205084
rect 480 204132 259520 204684
rect 560 203732 259520 204132
rect 480 201004 259520 203732
rect 480 200604 259440 201004
rect 480 199508 259520 200604
rect 560 199108 259520 199508
rect 480 196924 259520 199108
rect 480 196524 259440 196924
rect 480 194884 259520 196524
rect 560 194484 259520 194884
rect 480 192844 259520 194484
rect 480 192444 259440 192844
rect 480 190260 259520 192444
rect 560 189860 259520 190260
rect 480 188764 259520 189860
rect 480 188364 259440 188764
rect 480 185636 259520 188364
rect 560 185236 259520 185636
rect 480 184684 259520 185236
rect 480 184284 259440 184684
rect 480 181012 259520 184284
rect 560 180612 259520 181012
rect 480 180604 259520 180612
rect 480 180204 259440 180604
rect 480 176524 259520 180204
rect 480 176388 259440 176524
rect 560 176124 259440 176388
rect 560 175988 259520 176124
rect 480 172444 259520 175988
rect 480 172044 259440 172444
rect 480 171764 259520 172044
rect 560 171364 259520 171764
rect 480 168364 259520 171364
rect 480 167964 259440 168364
rect 480 167140 259520 167964
rect 560 166740 259520 167140
rect 480 164284 259520 166740
rect 480 163884 259440 164284
rect 480 162516 259520 163884
rect 560 162116 259520 162516
rect 480 160204 259520 162116
rect 480 159804 259440 160204
rect 480 157892 259520 159804
rect 560 157492 259520 157892
rect 480 156124 259520 157492
rect 480 155724 259440 156124
rect 480 153268 259520 155724
rect 560 152868 259520 153268
rect 480 152044 259520 152868
rect 480 151644 259440 152044
rect 480 148644 259520 151644
rect 560 148244 259520 148644
rect 480 147964 259520 148244
rect 480 147564 259440 147964
rect 480 144020 259520 147564
rect 560 143884 259520 144020
rect 560 143620 259440 143884
rect 480 143484 259440 143620
rect 480 139804 259520 143484
rect 480 139404 259440 139804
rect 480 139396 259520 139404
rect 560 138996 259520 139396
rect 480 135724 259520 138996
rect 480 135324 259440 135724
rect 480 134772 259520 135324
rect 560 134372 259520 134772
rect 480 131644 259520 134372
rect 480 131244 259440 131644
rect 480 130148 259520 131244
rect 560 129748 259520 130148
rect 480 127564 259520 129748
rect 480 127164 259440 127564
rect 480 125524 259520 127164
rect 560 125124 259520 125524
rect 480 123484 259520 125124
rect 480 123084 259440 123484
rect 480 120900 259520 123084
rect 560 120500 259520 120900
rect 480 119404 259520 120500
rect 480 119004 259440 119404
rect 480 116276 259520 119004
rect 560 115876 259520 116276
rect 480 115324 259520 115876
rect 480 114924 259440 115324
rect 480 111652 259520 114924
rect 560 111252 259520 111652
rect 480 111244 259520 111252
rect 480 110844 259440 111244
rect 480 107164 259520 110844
rect 480 107028 259440 107164
rect 560 106764 259440 107028
rect 560 106628 259520 106764
rect 480 103084 259520 106628
rect 480 102684 259440 103084
rect 480 102404 259520 102684
rect 560 102004 259520 102404
rect 480 99004 259520 102004
rect 480 98604 259440 99004
rect 480 97780 259520 98604
rect 560 97380 259520 97780
rect 480 94924 259520 97380
rect 480 94524 259440 94924
rect 480 93156 259520 94524
rect 560 92756 259520 93156
rect 480 90844 259520 92756
rect 480 90444 259440 90844
rect 480 88532 259520 90444
rect 560 88132 259520 88532
rect 480 86764 259520 88132
rect 480 86364 259440 86764
rect 480 83908 259520 86364
rect 560 83508 259520 83908
rect 480 82684 259520 83508
rect 480 82284 259440 82684
rect 480 79284 259520 82284
rect 560 78884 259520 79284
rect 480 78604 259520 78884
rect 480 78204 259440 78604
rect 480 74660 259520 78204
rect 560 74524 259520 74660
rect 560 74260 259440 74524
rect 480 74124 259440 74260
rect 480 70444 259520 74124
rect 480 70044 259440 70444
rect 480 70036 259520 70044
rect 560 69636 259520 70036
rect 480 66364 259520 69636
rect 480 65964 259440 66364
rect 480 65412 259520 65964
rect 560 65012 259520 65412
rect 480 62284 259520 65012
rect 480 61884 259440 62284
rect 480 60788 259520 61884
rect 560 60388 259520 60788
rect 480 58204 259520 60388
rect 480 57804 259440 58204
rect 480 56164 259520 57804
rect 560 55764 259520 56164
rect 480 54124 259520 55764
rect 480 53724 259440 54124
rect 480 51540 259520 53724
rect 560 51140 259520 51540
rect 480 50044 259520 51140
rect 480 49644 259440 50044
rect 480 46916 259520 49644
rect 560 46516 259520 46916
rect 480 45964 259520 46516
rect 480 45564 259440 45964
rect 480 42292 259520 45564
rect 560 41892 259520 42292
rect 480 41884 259520 41892
rect 480 41484 259440 41884
rect 480 37804 259520 41484
rect 480 37668 259440 37804
rect 560 37404 259440 37668
rect 560 37268 259520 37404
rect 480 33724 259520 37268
rect 480 33324 259440 33724
rect 480 33044 259520 33324
rect 560 32644 259520 33044
rect 480 29644 259520 32644
rect 480 29244 259440 29644
rect 480 28420 259520 29244
rect 560 28020 259520 28420
rect 480 25564 259520 28020
rect 480 25164 259440 25564
rect 480 23796 259520 25164
rect 560 23396 259520 23796
rect 480 21484 259520 23396
rect 480 21084 259440 21484
rect 480 19172 259520 21084
rect 560 18772 259520 19172
rect 480 17404 259520 18772
rect 480 17004 259440 17404
rect 480 14548 259520 17004
rect 560 14148 259520 14548
rect 480 13324 259520 14148
rect 480 12924 259440 13324
rect 480 9924 259520 12924
rect 560 9524 259520 9924
rect 480 9244 259520 9524
rect 480 8844 259440 9244
rect 480 5300 259520 8844
rect 560 5164 259520 5300
rect 560 4900 259440 5164
rect 480 4764 259440 4900
rect 480 2143 259520 4764
<< metal4 >>
rect 1794 2128 2414 317744
rect 7794 2128 8414 317744
rect 13794 2128 14414 317744
rect 19794 2128 20414 317744
rect 25794 2128 26414 317744
rect 31794 2128 32414 317744
rect 37794 2128 38414 317744
rect 43794 2128 44414 317744
rect 49794 2128 50414 317744
rect 55794 2128 56414 317744
rect 61794 2128 62414 317744
rect 67794 2128 68414 317744
rect 73794 2128 74414 317744
rect 79794 2128 80414 317744
rect 85794 2128 86414 317744
rect 91794 2128 92414 317744
rect 97794 2128 98414 317744
rect 103794 2128 104414 317744
rect 109794 2128 110414 317744
rect 115794 2128 116414 317744
rect 121794 2128 122414 317744
rect 127794 2128 128414 317744
rect 133794 2128 134414 317744
rect 139794 2128 140414 317744
rect 145794 2128 146414 317744
rect 151794 2128 152414 317744
rect 157794 2128 158414 317744
rect 163794 2128 164414 317744
rect 169794 2128 170414 317744
rect 175794 2128 176414 317744
rect 181794 2128 182414 317744
rect 187794 2128 188414 317744
rect 193794 2128 194414 317744
rect 199794 2128 200414 317744
rect 205794 2128 206414 317744
rect 211794 2128 212414 317744
rect 217794 2128 218414 317744
rect 223794 2128 224414 317744
rect 229794 2128 230414 317744
rect 235794 2128 236414 317744
rect 241794 2128 242414 317744
rect 247794 2128 248414 317744
rect 253794 2128 254414 317744
<< obsm4 >>
rect 97027 43283 97461 67693
<< labels >>
rlabel metal4 s 7794 2128 8414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 19794 2128 20414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 31794 2128 32414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 43794 2128 44414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67794 2128 68414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 79794 2128 80414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 103794 2128 104414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115794 2128 116414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127794 2128 128414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 139794 2128 140414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 151794 2128 152414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 163794 2128 164414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 175794 2128 176414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 187794 2128 188414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 199794 2128 200414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 211794 2128 212414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 223794 2128 224414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 235794 2128 236414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 247794 2128 248414 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13794 2128 14414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25794 2128 26414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 49794 2128 50414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 61794 2128 62414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 85794 2128 86414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 97794 2128 98414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 121794 2128 122414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 133794 2128 134414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145794 2128 146414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157794 2128 158414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 169794 2128 170414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 181794 2128 182414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 193794 2128 194414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 205794 2128 206414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217794 2128 218414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229794 2128 230414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 241794 2128 242414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 253794 2128 254414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 259520 135404 260960 135644 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 259520 257804 260960 258044 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 259520 270044 260960 270284 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 259520 282284 260960 282524 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 259520 294524 260960 294764 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 259520 306764 260960 307004 6 io_in[14]
port 8 nsew signal input
rlabel metal2 s 254278 319520 254390 320960 6 io_in[15]
port 9 nsew signal input
rlabel metal2 s 225574 319520 225686 320960 6 io_in[16]
port 10 nsew signal input
rlabel metal2 s 196870 319520 196982 320960 6 io_in[17]
port 11 nsew signal input
rlabel metal2 s 168166 319520 168278 320960 6 io_in[18]
port 12 nsew signal input
rlabel metal2 s 139462 319520 139574 320960 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 259520 147644 260960 147884 6 io_in[1]
port 14 nsew signal input
rlabel metal2 s 110758 319520 110870 320960 6 io_in[20]
port 15 nsew signal input
rlabel metal2 s 82054 319520 82166 320960 6 io_in[21]
port 16 nsew signal input
rlabel metal2 s 53350 319520 53462 320960 6 io_in[22]
port 17 nsew signal input
rlabel metal2 s 24646 319520 24758 320960 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s -960 314788 480 315028 4 io_in[24]
port 19 nsew signal input
rlabel metal3 s -960 300916 480 301156 4 io_in[25]
port 20 nsew signal input
rlabel metal3 s -960 287044 480 287284 4 io_in[26]
port 21 nsew signal input
rlabel metal3 s -960 273172 480 273412 4 io_in[27]
port 22 nsew signal input
rlabel metal3 s -960 259300 480 259540 4 io_in[28]
port 23 nsew signal input
rlabel metal3 s -960 245428 480 245668 4 io_in[29]
port 24 nsew signal input
rlabel metal3 s 259520 159884 260960 160124 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s -960 231556 480 231796 4 io_in[30]
port 26 nsew signal input
rlabel metal3 s -960 217684 480 217924 4 io_in[31]
port 27 nsew signal input
rlabel metal3 s -960 203812 480 204052 4 io_in[32]
port 28 nsew signal input
rlabel metal3 s -960 189940 480 190180 4 io_in[33]
port 29 nsew signal input
rlabel metal3 s -960 176068 480 176308 4 io_in[34]
port 30 nsew signal input
rlabel metal3 s -960 162196 480 162436 4 io_in[35]
port 31 nsew signal input
rlabel metal3 s 259520 172124 260960 172364 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 259520 184364 260960 184604 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 259520 196604 260960 196844 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 259520 208844 260960 209084 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 259520 221084 260960 221324 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 259520 233324 260960 233564 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 259520 245564 260960 245804 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 259520 143564 260960 143804 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 259520 265964 260960 266204 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 259520 278204 260960 278444 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 259520 290444 260960 290684 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 259520 302684 260960 302924 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 259520 314924 260960 315164 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 235142 319520 235254 320960 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 206438 319520 206550 320960 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 177734 319520 177846 320960 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 149030 319520 149142 320960 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 120326 319520 120438 320960 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 259520 155804 260960 156044 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 91622 319520 91734 320960 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 62918 319520 63030 320960 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 34214 319520 34326 320960 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5510 319520 5622 320960 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -960 305540 480 305780 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -960 291668 480 291908 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -960 277796 480 278036 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -960 263924 480 264164 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -960 250052 480 250292 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -960 236180 480 236420 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 259520 168044 260960 168284 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -960 222308 480 222548 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -960 208436 480 208676 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -960 194564 480 194804 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -960 180692 480 180932 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -960 166820 480 167060 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -960 152948 480 153188 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 259520 180284 260960 180524 6 io_oeb[3]
port 68 nsew signal output
rlabel metal3 s 259520 192524 260960 192764 6 io_oeb[4]
port 69 nsew signal output
rlabel metal3 s 259520 204764 260960 205004 6 io_oeb[5]
port 70 nsew signal output
rlabel metal3 s 259520 217004 260960 217244 6 io_oeb[6]
port 71 nsew signal output
rlabel metal3 s 259520 229244 260960 229484 6 io_oeb[7]
port 72 nsew signal output
rlabel metal3 s 259520 241484 260960 241724 6 io_oeb[8]
port 73 nsew signal output
rlabel metal3 s 259520 253724 260960 253964 6 io_oeb[9]
port 74 nsew signal output
rlabel metal3 s 259520 139484 260960 139724 6 io_out[0]
port 75 nsew signal output
rlabel metal3 s 259520 261884 260960 262124 6 io_out[10]
port 76 nsew signal output
rlabel metal3 s 259520 274124 260960 274364 6 io_out[11]
port 77 nsew signal output
rlabel metal3 s 259520 286364 260960 286604 6 io_out[12]
port 78 nsew signal output
rlabel metal3 s 259520 298604 260960 298844 6 io_out[13]
port 79 nsew signal output
rlabel metal3 s 259520 310844 260960 311084 6 io_out[14]
port 80 nsew signal output
rlabel metal2 s 244710 319520 244822 320960 6 io_out[15]
port 81 nsew signal output
rlabel metal2 s 216006 319520 216118 320960 6 io_out[16]
port 82 nsew signal output
rlabel metal2 s 187302 319520 187414 320960 6 io_out[17]
port 83 nsew signal output
rlabel metal2 s 158598 319520 158710 320960 6 io_out[18]
port 84 nsew signal output
rlabel metal2 s 129894 319520 130006 320960 6 io_out[19]
port 85 nsew signal output
rlabel metal3 s 259520 151724 260960 151964 6 io_out[1]
port 86 nsew signal output
rlabel metal2 s 101190 319520 101302 320960 6 io_out[20]
port 87 nsew signal output
rlabel metal2 s 72486 319520 72598 320960 6 io_out[21]
port 88 nsew signal output
rlabel metal2 s 43782 319520 43894 320960 6 io_out[22]
port 89 nsew signal output
rlabel metal2 s 15078 319520 15190 320960 6 io_out[23]
port 90 nsew signal output
rlabel metal3 s -960 310164 480 310404 4 io_out[24]
port 91 nsew signal output
rlabel metal3 s -960 296292 480 296532 4 io_out[25]
port 92 nsew signal output
rlabel metal3 s -960 282420 480 282660 4 io_out[26]
port 93 nsew signal output
rlabel metal3 s -960 268548 480 268788 4 io_out[27]
port 94 nsew signal output
rlabel metal3 s -960 254676 480 254916 4 io_out[28]
port 95 nsew signal output
rlabel metal3 s -960 240804 480 241044 4 io_out[29]
port 96 nsew signal output
rlabel metal3 s 259520 163964 260960 164204 6 io_out[2]
port 97 nsew signal output
rlabel metal3 s -960 226932 480 227172 4 io_out[30]
port 98 nsew signal output
rlabel metal3 s -960 213060 480 213300 4 io_out[31]
port 99 nsew signal output
rlabel metal3 s -960 199188 480 199428 4 io_out[32]
port 100 nsew signal output
rlabel metal3 s -960 185316 480 185556 4 io_out[33]
port 101 nsew signal output
rlabel metal3 s -960 171444 480 171684 4 io_out[34]
port 102 nsew signal output
rlabel metal3 s -960 157572 480 157812 4 io_out[35]
port 103 nsew signal output
rlabel metal3 s 259520 176204 260960 176444 6 io_out[3]
port 104 nsew signal output
rlabel metal3 s 259520 188444 260960 188684 6 io_out[4]
port 105 nsew signal output
rlabel metal3 s 259520 200684 260960 200924 6 io_out[5]
port 106 nsew signal output
rlabel metal3 s 259520 212924 260960 213164 6 io_out[6]
port 107 nsew signal output
rlabel metal3 s 259520 225164 260960 225404 6 io_out[7]
port 108 nsew signal output
rlabel metal3 s 259520 237404 260960 237644 6 io_out[8]
port 109 nsew signal output
rlabel metal3 s 259520 249644 260960 249884 6 io_out[9]
port 110 nsew signal output
rlabel metal3 s -960 148324 480 148564 4 la_data_in[0]
port 111 nsew signal input
rlabel metal3 s -960 102084 480 102324 4 la_data_in[10]
port 112 nsew signal input
rlabel metal3 s -960 97460 480 97700 4 la_data_in[11]
port 113 nsew signal input
rlabel metal3 s -960 92836 480 93076 4 la_data_in[12]
port 114 nsew signal input
rlabel metal3 s -960 88212 480 88452 4 la_data_in[13]
port 115 nsew signal input
rlabel metal3 s -960 83588 480 83828 4 la_data_in[14]
port 116 nsew signal input
rlabel metal3 s -960 78964 480 79204 4 la_data_in[15]
port 117 nsew signal input
rlabel metal3 s -960 74340 480 74580 4 la_data_in[16]
port 118 nsew signal input
rlabel metal3 s -960 69716 480 69956 4 la_data_in[17]
port 119 nsew signal input
rlabel metal3 s -960 65092 480 65332 4 la_data_in[18]
port 120 nsew signal input
rlabel metal3 s -960 60468 480 60708 4 la_data_in[19]
port 121 nsew signal input
rlabel metal3 s -960 143700 480 143940 4 la_data_in[1]
port 122 nsew signal input
rlabel metal3 s -960 55844 480 56084 4 la_data_in[20]
port 123 nsew signal input
rlabel metal3 s -960 51220 480 51460 4 la_data_in[21]
port 124 nsew signal input
rlabel metal3 s -960 46596 480 46836 4 la_data_in[22]
port 125 nsew signal input
rlabel metal3 s -960 41972 480 42212 4 la_data_in[23]
port 126 nsew signal input
rlabel metal3 s -960 37348 480 37588 4 la_data_in[24]
port 127 nsew signal input
rlabel metal3 s -960 32724 480 32964 4 la_data_in[25]
port 128 nsew signal input
rlabel metal3 s -960 28100 480 28340 4 la_data_in[26]
port 129 nsew signal input
rlabel metal3 s -960 23476 480 23716 4 la_data_in[27]
port 130 nsew signal input
rlabel metal3 s -960 18852 480 19092 4 la_data_in[28]
port 131 nsew signal input
rlabel metal3 s -960 14228 480 14468 4 la_data_in[29]
port 132 nsew signal input
rlabel metal3 s -960 139076 480 139316 4 la_data_in[2]
port 133 nsew signal input
rlabel metal3 s -960 9604 480 9844 4 la_data_in[30]
port 134 nsew signal input
rlabel metal3 s -960 4980 480 5220 4 la_data_in[31]
port 135 nsew signal input
rlabel metal3 s -960 134452 480 134692 4 la_data_in[3]
port 136 nsew signal input
rlabel metal3 s -960 129828 480 130068 4 la_data_in[4]
port 137 nsew signal input
rlabel metal3 s -960 125204 480 125444 4 la_data_in[5]
port 138 nsew signal input
rlabel metal3 s -960 120580 480 120820 4 la_data_in[6]
port 139 nsew signal input
rlabel metal3 s -960 115956 480 116196 4 la_data_in[7]
port 140 nsew signal input
rlabel metal3 s -960 111332 480 111572 4 la_data_in[8]
port 141 nsew signal input
rlabel metal3 s -960 106708 480 106948 4 la_data_in[9]
port 142 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[0]
port 143 nsew signal output
rlabel metal2 s 209474 -960 209586 480 8 la_data_out[10]
port 144 nsew signal output
rlabel metal2 s 211222 -960 211334 480 8 la_data_out[11]
port 145 nsew signal output
rlabel metal2 s 212970 -960 213082 480 8 la_data_out[12]
port 146 nsew signal output
rlabel metal2 s 214718 -960 214830 480 8 la_data_out[13]
port 147 nsew signal output
rlabel metal2 s 216466 -960 216578 480 8 la_data_out[14]
port 148 nsew signal output
rlabel metal2 s 218214 -960 218326 480 8 la_data_out[15]
port 149 nsew signal output
rlabel metal2 s 219962 -960 220074 480 8 la_data_out[16]
port 150 nsew signal output
rlabel metal2 s 221710 -960 221822 480 8 la_data_out[17]
port 151 nsew signal output
rlabel metal2 s 223458 -960 223570 480 8 la_data_out[18]
port 152 nsew signal output
rlabel metal2 s 225206 -960 225318 480 8 la_data_out[19]
port 153 nsew signal output
rlabel metal2 s 193742 -960 193854 480 8 la_data_out[1]
port 154 nsew signal output
rlabel metal2 s 226954 -960 227066 480 8 la_data_out[20]
port 155 nsew signal output
rlabel metal2 s 228702 -960 228814 480 8 la_data_out[21]
port 156 nsew signal output
rlabel metal2 s 230450 -960 230562 480 8 la_data_out[22]
port 157 nsew signal output
rlabel metal2 s 232198 -960 232310 480 8 la_data_out[23]
port 158 nsew signal output
rlabel metal2 s 233946 -960 234058 480 8 la_data_out[24]
port 159 nsew signal output
rlabel metal2 s 235694 -960 235806 480 8 la_data_out[25]
port 160 nsew signal output
rlabel metal2 s 237442 -960 237554 480 8 la_data_out[26]
port 161 nsew signal output
rlabel metal2 s 239190 -960 239302 480 8 la_data_out[27]
port 162 nsew signal output
rlabel metal2 s 240938 -960 241050 480 8 la_data_out[28]
port 163 nsew signal output
rlabel metal2 s 242686 -960 242798 480 8 la_data_out[29]
port 164 nsew signal output
rlabel metal2 s 195490 -960 195602 480 8 la_data_out[2]
port 165 nsew signal output
rlabel metal2 s 244434 -960 244546 480 8 la_data_out[30]
port 166 nsew signal output
rlabel metal2 s 246182 -960 246294 480 8 la_data_out[31]
port 167 nsew signal output
rlabel metal2 s 197238 -960 197350 480 8 la_data_out[3]
port 168 nsew signal output
rlabel metal2 s 198986 -960 199098 480 8 la_data_out[4]
port 169 nsew signal output
rlabel metal2 s 200734 -960 200846 480 8 la_data_out[5]
port 170 nsew signal output
rlabel metal2 s 202482 -960 202594 480 8 la_data_out[6]
port 171 nsew signal output
rlabel metal2 s 204230 -960 204342 480 8 la_data_out[7]
port 172 nsew signal output
rlabel metal2 s 205978 -960 206090 480 8 la_data_out[8]
port 173 nsew signal output
rlabel metal2 s 207726 -960 207838 480 8 la_data_out[9]
port 174 nsew signal output
rlabel metal3 s 259520 4844 260960 5084 6 la_oenb[0]
port 175 nsew signal input
rlabel metal3 s 259520 45644 260960 45884 6 la_oenb[10]
port 176 nsew signal input
rlabel metal3 s 259520 49724 260960 49964 6 la_oenb[11]
port 177 nsew signal input
rlabel metal3 s 259520 53804 260960 54044 6 la_oenb[12]
port 178 nsew signal input
rlabel metal3 s 259520 57884 260960 58124 6 la_oenb[13]
port 179 nsew signal input
rlabel metal3 s 259520 61964 260960 62204 6 la_oenb[14]
port 180 nsew signal input
rlabel metal3 s 259520 66044 260960 66284 6 la_oenb[15]
port 181 nsew signal input
rlabel metal3 s 259520 70124 260960 70364 6 la_oenb[16]
port 182 nsew signal input
rlabel metal3 s 259520 74204 260960 74444 6 la_oenb[17]
port 183 nsew signal input
rlabel metal3 s 259520 78284 260960 78524 6 la_oenb[18]
port 184 nsew signal input
rlabel metal3 s 259520 82364 260960 82604 6 la_oenb[19]
port 185 nsew signal input
rlabel metal3 s 259520 8924 260960 9164 6 la_oenb[1]
port 186 nsew signal input
rlabel metal3 s 259520 86444 260960 86684 6 la_oenb[20]
port 187 nsew signal input
rlabel metal3 s 259520 90524 260960 90764 6 la_oenb[21]
port 188 nsew signal input
rlabel metal3 s 259520 94604 260960 94844 6 la_oenb[22]
port 189 nsew signal input
rlabel metal3 s 259520 98684 260960 98924 6 la_oenb[23]
port 190 nsew signal input
rlabel metal3 s 259520 102764 260960 103004 6 la_oenb[24]
port 191 nsew signal input
rlabel metal3 s 259520 106844 260960 107084 6 la_oenb[25]
port 192 nsew signal input
rlabel metal3 s 259520 110924 260960 111164 6 la_oenb[26]
port 193 nsew signal input
rlabel metal3 s 259520 115004 260960 115244 6 la_oenb[27]
port 194 nsew signal input
rlabel metal3 s 259520 119084 260960 119324 6 la_oenb[28]
port 195 nsew signal input
rlabel metal3 s 259520 123164 260960 123404 6 la_oenb[29]
port 196 nsew signal input
rlabel metal3 s 259520 13004 260960 13244 6 la_oenb[2]
port 197 nsew signal input
rlabel metal3 s 259520 127244 260960 127484 6 la_oenb[30]
port 198 nsew signal input
rlabel metal3 s 259520 131324 260960 131564 6 la_oenb[31]
port 199 nsew signal input
rlabel metal3 s 259520 17084 260960 17324 6 la_oenb[3]
port 200 nsew signal input
rlabel metal3 s 259520 21164 260960 21404 6 la_oenb[4]
port 201 nsew signal input
rlabel metal3 s 259520 25244 260960 25484 6 la_oenb[5]
port 202 nsew signal input
rlabel metal3 s 259520 29324 260960 29564 6 la_oenb[6]
port 203 nsew signal input
rlabel metal3 s 259520 33404 260960 33644 6 la_oenb[7]
port 204 nsew signal input
rlabel metal3 s 259520 37484 260960 37724 6 la_oenb[8]
port 205 nsew signal input
rlabel metal3 s 259520 41564 260960 41804 6 la_oenb[9]
port 206 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 user_clock2
port 207 nsew signal input
rlabel metal2 s 249678 -960 249790 480 8 user_irq[0]
port 208 nsew signal output
rlabel metal2 s 251426 -960 251538 480 8 user_irq[1]
port 209 nsew signal output
rlabel metal2 s 253174 -960 253286 480 8 user_irq[2]
port 210 nsew signal output
rlabel metal2 s 6706 -960 6818 480 8 wb_clk_i
port 211 nsew signal input
rlabel metal2 s 8454 -960 8566 480 8 wb_rst_i
port 212 nsew signal input
rlabel metal2 s 10202 -960 10314 480 8 wbs_ack_o
port 213 nsew signal output
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[0]
port 214 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[10]
port 215 nsew signal input
rlabel metal2 s 81870 -960 81982 480 8 wbs_adr_i[11]
port 216 nsew signal input
rlabel metal2 s 87114 -960 87226 480 8 wbs_adr_i[12]
port 217 nsew signal input
rlabel metal2 s 92358 -960 92470 480 8 wbs_adr_i[13]
port 218 nsew signal input
rlabel metal2 s 97602 -960 97714 480 8 wbs_adr_i[14]
port 219 nsew signal input
rlabel metal2 s 102846 -960 102958 480 8 wbs_adr_i[15]
port 220 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[16]
port 221 nsew signal input
rlabel metal2 s 113334 -960 113446 480 8 wbs_adr_i[17]
port 222 nsew signal input
rlabel metal2 s 118578 -960 118690 480 8 wbs_adr_i[18]
port 223 nsew signal input
rlabel metal2 s 123822 -960 123934 480 8 wbs_adr_i[19]
port 224 nsew signal input
rlabel metal2 s 24186 -960 24298 480 8 wbs_adr_i[1]
port 225 nsew signal input
rlabel metal2 s 129066 -960 129178 480 8 wbs_adr_i[20]
port 226 nsew signal input
rlabel metal2 s 134310 -960 134422 480 8 wbs_adr_i[21]
port 227 nsew signal input
rlabel metal2 s 139554 -960 139666 480 8 wbs_adr_i[22]
port 228 nsew signal input
rlabel metal2 s 144798 -960 144910 480 8 wbs_adr_i[23]
port 229 nsew signal input
rlabel metal2 s 150042 -960 150154 480 8 wbs_adr_i[24]
port 230 nsew signal input
rlabel metal2 s 155286 -960 155398 480 8 wbs_adr_i[25]
port 231 nsew signal input
rlabel metal2 s 160530 -960 160642 480 8 wbs_adr_i[26]
port 232 nsew signal input
rlabel metal2 s 165774 -960 165886 480 8 wbs_adr_i[27]
port 233 nsew signal input
rlabel metal2 s 171018 -960 171130 480 8 wbs_adr_i[28]
port 234 nsew signal input
rlabel metal2 s 176262 -960 176374 480 8 wbs_adr_i[29]
port 235 nsew signal input
rlabel metal2 s 31178 -960 31290 480 8 wbs_adr_i[2]
port 236 nsew signal input
rlabel metal2 s 181506 -960 181618 480 8 wbs_adr_i[30]
port 237 nsew signal input
rlabel metal2 s 186750 -960 186862 480 8 wbs_adr_i[31]
port 238 nsew signal input
rlabel metal2 s 38170 -960 38282 480 8 wbs_adr_i[3]
port 239 nsew signal input
rlabel metal2 s 45162 -960 45274 480 8 wbs_adr_i[4]
port 240 nsew signal input
rlabel metal2 s 50406 -960 50518 480 8 wbs_adr_i[5]
port 241 nsew signal input
rlabel metal2 s 55650 -960 55762 480 8 wbs_adr_i[6]
port 242 nsew signal input
rlabel metal2 s 60894 -960 61006 480 8 wbs_adr_i[7]
port 243 nsew signal input
rlabel metal2 s 66138 -960 66250 480 8 wbs_adr_i[8]
port 244 nsew signal input
rlabel metal2 s 71382 -960 71494 480 8 wbs_adr_i[9]
port 245 nsew signal input
rlabel metal2 s 11950 -960 12062 480 8 wbs_cyc_i
port 246 nsew signal input
rlabel metal2 s 18942 -960 19054 480 8 wbs_dat_i[0]
port 247 nsew signal input
rlabel metal2 s 78374 -960 78486 480 8 wbs_dat_i[10]
port 248 nsew signal input
rlabel metal2 s 83618 -960 83730 480 8 wbs_dat_i[11]
port 249 nsew signal input
rlabel metal2 s 88862 -960 88974 480 8 wbs_dat_i[12]
port 250 nsew signal input
rlabel metal2 s 94106 -960 94218 480 8 wbs_dat_i[13]
port 251 nsew signal input
rlabel metal2 s 99350 -960 99462 480 8 wbs_dat_i[14]
port 252 nsew signal input
rlabel metal2 s 104594 -960 104706 480 8 wbs_dat_i[15]
port 253 nsew signal input
rlabel metal2 s 109838 -960 109950 480 8 wbs_dat_i[16]
port 254 nsew signal input
rlabel metal2 s 115082 -960 115194 480 8 wbs_dat_i[17]
port 255 nsew signal input
rlabel metal2 s 120326 -960 120438 480 8 wbs_dat_i[18]
port 256 nsew signal input
rlabel metal2 s 125570 -960 125682 480 8 wbs_dat_i[19]
port 257 nsew signal input
rlabel metal2 s 25934 -960 26046 480 8 wbs_dat_i[1]
port 258 nsew signal input
rlabel metal2 s 130814 -960 130926 480 8 wbs_dat_i[20]
port 259 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 wbs_dat_i[21]
port 260 nsew signal input
rlabel metal2 s 141302 -960 141414 480 8 wbs_dat_i[22]
port 261 nsew signal input
rlabel metal2 s 146546 -960 146658 480 8 wbs_dat_i[23]
port 262 nsew signal input
rlabel metal2 s 151790 -960 151902 480 8 wbs_dat_i[24]
port 263 nsew signal input
rlabel metal2 s 157034 -960 157146 480 8 wbs_dat_i[25]
port 264 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 wbs_dat_i[26]
port 265 nsew signal input
rlabel metal2 s 167522 -960 167634 480 8 wbs_dat_i[27]
port 266 nsew signal input
rlabel metal2 s 172766 -960 172878 480 8 wbs_dat_i[28]
port 267 nsew signal input
rlabel metal2 s 178010 -960 178122 480 8 wbs_dat_i[29]
port 268 nsew signal input
rlabel metal2 s 32926 -960 33038 480 8 wbs_dat_i[2]
port 269 nsew signal input
rlabel metal2 s 183254 -960 183366 480 8 wbs_dat_i[30]
port 270 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 wbs_dat_i[31]
port 271 nsew signal input
rlabel metal2 s 39918 -960 40030 480 8 wbs_dat_i[3]
port 272 nsew signal input
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_i[4]
port 273 nsew signal input
rlabel metal2 s 52154 -960 52266 480 8 wbs_dat_i[5]
port 274 nsew signal input
rlabel metal2 s 57398 -960 57510 480 8 wbs_dat_i[6]
port 275 nsew signal input
rlabel metal2 s 62642 -960 62754 480 8 wbs_dat_i[7]
port 276 nsew signal input
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_i[8]
port 277 nsew signal input
rlabel metal2 s 73130 -960 73242 480 8 wbs_dat_i[9]
port 278 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_dat_o[0]
port 279 nsew signal output
rlabel metal2 s 80122 -960 80234 480 8 wbs_dat_o[10]
port 280 nsew signal output
rlabel metal2 s 85366 -960 85478 480 8 wbs_dat_o[11]
port 281 nsew signal output
rlabel metal2 s 90610 -960 90722 480 8 wbs_dat_o[12]
port 282 nsew signal output
rlabel metal2 s 95854 -960 95966 480 8 wbs_dat_o[13]
port 283 nsew signal output
rlabel metal2 s 101098 -960 101210 480 8 wbs_dat_o[14]
port 284 nsew signal output
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_o[15]
port 285 nsew signal output
rlabel metal2 s 111586 -960 111698 480 8 wbs_dat_o[16]
port 286 nsew signal output
rlabel metal2 s 116830 -960 116942 480 8 wbs_dat_o[17]
port 287 nsew signal output
rlabel metal2 s 122074 -960 122186 480 8 wbs_dat_o[18]
port 288 nsew signal output
rlabel metal2 s 127318 -960 127430 480 8 wbs_dat_o[19]
port 289 nsew signal output
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_o[1]
port 290 nsew signal output
rlabel metal2 s 132562 -960 132674 480 8 wbs_dat_o[20]
port 291 nsew signal output
rlabel metal2 s 137806 -960 137918 480 8 wbs_dat_o[21]
port 292 nsew signal output
rlabel metal2 s 143050 -960 143162 480 8 wbs_dat_o[22]
port 293 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 wbs_dat_o[23]
port 294 nsew signal output
rlabel metal2 s 153538 -960 153650 480 8 wbs_dat_o[24]
port 295 nsew signal output
rlabel metal2 s 158782 -960 158894 480 8 wbs_dat_o[25]
port 296 nsew signal output
rlabel metal2 s 164026 -960 164138 480 8 wbs_dat_o[26]
port 297 nsew signal output
rlabel metal2 s 169270 -960 169382 480 8 wbs_dat_o[27]
port 298 nsew signal output
rlabel metal2 s 174514 -960 174626 480 8 wbs_dat_o[28]
port 299 nsew signal output
rlabel metal2 s 179758 -960 179870 480 8 wbs_dat_o[29]
port 300 nsew signal output
rlabel metal2 s 34674 -960 34786 480 8 wbs_dat_o[2]
port 301 nsew signal output
rlabel metal2 s 185002 -960 185114 480 8 wbs_dat_o[30]
port 302 nsew signal output
rlabel metal2 s 190246 -960 190358 480 8 wbs_dat_o[31]
port 303 nsew signal output
rlabel metal2 s 41666 -960 41778 480 8 wbs_dat_o[3]
port 304 nsew signal output
rlabel metal2 s 48658 -960 48770 480 8 wbs_dat_o[4]
port 305 nsew signal output
rlabel metal2 s 53902 -960 54014 480 8 wbs_dat_o[5]
port 306 nsew signal output
rlabel metal2 s 59146 -960 59258 480 8 wbs_dat_o[6]
port 307 nsew signal output
rlabel metal2 s 64390 -960 64502 480 8 wbs_dat_o[7]
port 308 nsew signal output
rlabel metal2 s 69634 -960 69746 480 8 wbs_dat_o[8]
port 309 nsew signal output
rlabel metal2 s 74878 -960 74990 480 8 wbs_dat_o[9]
port 310 nsew signal output
rlabel metal2 s 22438 -960 22550 480 8 wbs_sel_i[0]
port 311 nsew signal input
rlabel metal2 s 29430 -960 29542 480 8 wbs_sel_i[1]
port 312 nsew signal input
rlabel metal2 s 36422 -960 36534 480 8 wbs_sel_i[2]
port 313 nsew signal input
rlabel metal2 s 43414 -960 43526 480 8 wbs_sel_i[3]
port 314 nsew signal input
rlabel metal2 s 13698 -960 13810 480 8 wbs_stb_i
port 315 nsew signal input
rlabel metal2 s 15446 -960 15558 480 8 wbs_we_i
port 316 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 260000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 39787608
string GDS_FILE /home/hosni/mpc/openlane/user_project_5/runs/23_04_23_18_35/results/signoff/user_project_5.magic.gds
string GDS_START 453092
<< end >>

